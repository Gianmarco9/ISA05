`ifndef MY_DEFINES
	`define MY_DEFINES
		parameter nb=32;
		parameter n_prod=64;
`endif
