`ifndef MY_DEFINES
	`define MY_DEFINES
		parameter nb=32;
		parameter n_prod=32;
		parameter pipe_stages=6;
`endif
