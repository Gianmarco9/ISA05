LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE work.mypackage.all;

ENTITY dadda_tree IS
PORT(	PP_IN: IN DADDA_ARRAY;
	PP_OUT1:OUT STD_LOGIC_VECTOR(n_prod-1 DOWNTO 0);
	PP_OUT2:OUT STD_LOGIC_VECTOR(n_prod-1 DOWNTO 0)
);
END ENTITY;


ARCHITECTURE struct OF dadda_tree IS

COMPONENT FA 
PORT(	A: IN STD_LOGIC;
	B: IN STD_LOGIC;
	Ci: IN STD_LOGIC;
	S: OUT STD_LOGIC;
	Co: OUT STD_LOGIC);
END COMPONENT;
	
COMPONENT HA 
PORT(	A: IN STD_LOGIC;
	B: IN STD_LOGIC;
	S: OUT STD_LOGIC;
	Co: OUT STD_LOGIC);
END COMPONENT;

SIGNAL HA_lev6_col24_inst0_port_S: std_logic;
SIGNAL HA_lev6_col24_inst0_port_COUT: std_logic;
SIGNAL HA_lev6_col25_inst0_port_S: std_logic;
SIGNAL HA_lev6_col25_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col26_inst0_port_S: std_logic;
SIGNAL FA_lev6_col26_inst0_port_COUT: std_logic;
SIGNAL HA_lev6_col26_inst1_port_S: std_logic;
SIGNAL HA_lev6_col26_inst1_port_COUT: std_logic;
SIGNAL FA_lev6_col27_inst0_port_S: std_logic;
SIGNAL FA_lev6_col27_inst0_port_COUT: std_logic;
SIGNAL HA_lev6_col27_inst1_port_S: std_logic;
SIGNAL HA_lev6_col27_inst1_port_COUT: std_logic;
SIGNAL FA_lev6_col28_inst0_port_S: std_logic;
SIGNAL FA_lev6_col28_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col28_inst1_port_S: std_logic;
SIGNAL FA_lev6_col28_inst1_port_COUT: std_logic;
SIGNAL HA_lev6_col28_inst2_port_S: std_logic;
SIGNAL HA_lev6_col28_inst2_port_COUT: std_logic;
SIGNAL FA_lev6_col29_inst0_port_S: std_logic;
SIGNAL FA_lev6_col29_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col29_inst1_port_S: std_logic;
SIGNAL FA_lev6_col29_inst1_port_COUT: std_logic;
SIGNAL HA_lev6_col29_inst2_port_S: std_logic;
SIGNAL HA_lev6_col29_inst2_port_COUT: std_logic;
SIGNAL FA_lev6_col30_inst0_port_S: std_logic;
SIGNAL FA_lev6_col30_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col30_inst1_port_S: std_logic;
SIGNAL FA_lev6_col30_inst1_port_COUT: std_logic;
SIGNAL FA_lev6_col30_inst2_port_S: std_logic;
SIGNAL FA_lev6_col30_inst2_port_COUT: std_logic;
SIGNAL HA_lev6_col30_inst3_port_S: std_logic;
SIGNAL HA_lev6_col30_inst3_port_COUT: std_logic;
SIGNAL FA_lev6_col31_inst0_port_S: std_logic;
SIGNAL FA_lev6_col31_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col31_inst1_port_S: std_logic;
SIGNAL FA_lev6_col31_inst1_port_COUT: std_logic;
SIGNAL FA_lev6_col31_inst2_port_S: std_logic;
SIGNAL FA_lev6_col31_inst2_port_COUT: std_logic;
SIGNAL HA_lev6_col31_inst3_port_S: std_logic;
SIGNAL HA_lev6_col31_inst3_port_COUT: std_logic;
SIGNAL FA_lev6_col32_inst0_port_S: std_logic;
SIGNAL FA_lev6_col32_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col32_inst1_port_S: std_logic;
SIGNAL FA_lev6_col32_inst1_port_COUT: std_logic;
SIGNAL FA_lev6_col32_inst2_port_S: std_logic;
SIGNAL FA_lev6_col32_inst2_port_COUT: std_logic;
SIGNAL FA_lev6_col32_inst3_port_S: std_logic;
SIGNAL FA_lev6_col32_inst3_port_COUT: std_logic;
SIGNAL FA_lev6_col33_inst0_port_S: std_logic;
SIGNAL FA_lev6_col33_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col33_inst1_port_S: std_logic;
SIGNAL FA_lev6_col33_inst1_port_COUT: std_logic;
SIGNAL FA_lev6_col33_inst2_port_S: std_logic;
SIGNAL FA_lev6_col33_inst2_port_COUT: std_logic;
SIGNAL FA_lev6_col33_inst3_port_S: std_logic;
SIGNAL FA_lev6_col33_inst3_port_COUT: std_logic;
SIGNAL FA_lev6_col34_inst0_port_S: std_logic;
SIGNAL FA_lev6_col34_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col34_inst1_port_S: std_logic;
SIGNAL FA_lev6_col34_inst1_port_COUT: std_logic;
SIGNAL FA_lev6_col34_inst2_port_S: std_logic;
SIGNAL FA_lev6_col34_inst2_port_COUT: std_logic;
SIGNAL FA_lev6_col34_inst3_port_S: std_logic;
SIGNAL FA_lev6_col34_inst3_port_COUT: std_logic;
SIGNAL FA_lev6_col35_inst0_port_S: std_logic;
SIGNAL FA_lev6_col35_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col35_inst1_port_S: std_logic;
SIGNAL FA_lev6_col35_inst1_port_COUT: std_logic;
SIGNAL FA_lev6_col35_inst2_port_S: std_logic;
SIGNAL FA_lev6_col35_inst2_port_COUT: std_logic;
SIGNAL FA_lev6_col35_inst3_port_S: std_logic;
SIGNAL FA_lev6_col35_inst3_port_COUT: std_logic;
SIGNAL FA_lev6_col36_inst0_port_S: std_logic;
SIGNAL FA_lev6_col36_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col36_inst1_port_S: std_logic;
SIGNAL FA_lev6_col36_inst1_port_COUT: std_logic;
SIGNAL FA_lev6_col36_inst2_port_S: std_logic;
SIGNAL FA_lev6_col36_inst2_port_COUT: std_logic;
SIGNAL HA_lev6_col36_inst3_port_S: std_logic;
SIGNAL HA_lev6_col36_inst3_port_COUT: std_logic;
SIGNAL FA_lev6_col37_inst0_port_S: std_logic;
SIGNAL FA_lev6_col37_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col37_inst1_port_S: std_logic;
SIGNAL FA_lev6_col37_inst1_port_COUT: std_logic;
SIGNAL FA_lev6_col37_inst2_port_S: std_logic;
SIGNAL FA_lev6_col37_inst2_port_COUT: std_logic;
SIGNAL FA_lev6_col38_inst0_port_S: std_logic;
SIGNAL FA_lev6_col38_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col38_inst1_port_S: std_logic;
SIGNAL FA_lev6_col38_inst1_port_COUT: std_logic;
SIGNAL HA_lev6_col38_inst2_port_S: std_logic;
SIGNAL HA_lev6_col38_inst2_port_COUT: std_logic;
SIGNAL FA_lev6_col39_inst0_port_S: std_logic;
SIGNAL FA_lev6_col39_inst0_port_COUT: std_logic;
SIGNAL FA_lev6_col39_inst1_port_S: std_logic;
SIGNAL FA_lev6_col39_inst1_port_COUT: std_logic;
SIGNAL FA_lev6_col40_inst0_port_S: std_logic;
SIGNAL FA_lev6_col40_inst0_port_COUT: std_logic;
SIGNAL HA_lev6_col40_inst1_port_S: std_logic;
SIGNAL HA_lev6_col40_inst1_port_COUT: std_logic;
SIGNAL FA_lev6_col41_inst0_port_S: std_logic;
SIGNAL FA_lev6_col41_inst0_port_COUT: std_logic;
SIGNAL HA_lev6_col42_inst0_port_S: std_logic;
SIGNAL HA_lev6_col42_inst0_port_COUT: std_logic;
SIGNAL HA_lev5_col16_inst0_port_S: std_logic;
SIGNAL HA_lev5_col16_inst0_port_COUT: std_logic;
SIGNAL HA_lev5_col17_inst0_port_S: std_logic;
SIGNAL HA_lev5_col17_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col18_inst0_port_S: std_logic;
SIGNAL FA_lev5_col18_inst0_port_COUT: std_logic;
SIGNAL HA_lev5_col18_inst1_port_S: std_logic;
SIGNAL HA_lev5_col18_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col19_inst0_port_S: std_logic;
SIGNAL FA_lev5_col19_inst0_port_COUT: std_logic;
SIGNAL HA_lev5_col19_inst1_port_S: std_logic;
SIGNAL HA_lev5_col19_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col20_inst0_port_S: std_logic;
SIGNAL FA_lev5_col20_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col20_inst1_port_S: std_logic;
SIGNAL FA_lev5_col20_inst1_port_COUT: std_logic;
SIGNAL HA_lev5_col20_inst2_port_S: std_logic;
SIGNAL HA_lev5_col20_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col21_inst0_port_S: std_logic;
SIGNAL FA_lev5_col21_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col21_inst1_port_S: std_logic;
SIGNAL FA_lev5_col21_inst1_port_COUT: std_logic;
SIGNAL HA_lev5_col21_inst2_port_S: std_logic;
SIGNAL HA_lev5_col21_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col22_inst0_port_S: std_logic;
SIGNAL FA_lev5_col22_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col22_inst1_port_S: std_logic;
SIGNAL FA_lev5_col22_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col22_inst2_port_S: std_logic;
SIGNAL FA_lev5_col22_inst2_port_COUT: std_logic;
SIGNAL HA_lev5_col22_inst3_port_S: std_logic;
SIGNAL HA_lev5_col22_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col23_inst0_port_S: std_logic;
SIGNAL FA_lev5_col23_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col23_inst1_port_S: std_logic;
SIGNAL FA_lev5_col23_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col23_inst2_port_S: std_logic;
SIGNAL FA_lev5_col23_inst2_port_COUT: std_logic;
SIGNAL HA_lev5_col23_inst3_port_S: std_logic;
SIGNAL HA_lev5_col23_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col24_inst0_port_S: std_logic;
SIGNAL FA_lev5_col24_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col24_inst1_port_S: std_logic;
SIGNAL FA_lev5_col24_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col24_inst2_port_S: std_logic;
SIGNAL FA_lev5_col24_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col24_inst3_port_S: std_logic;
SIGNAL FA_lev5_col24_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col25_inst0_port_S: std_logic;
SIGNAL FA_lev5_col25_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col25_inst1_port_S: std_logic;
SIGNAL FA_lev5_col25_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col25_inst2_port_S: std_logic;
SIGNAL FA_lev5_col25_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col25_inst3_port_S: std_logic;
SIGNAL FA_lev5_col25_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col26_inst0_port_S: std_logic;
SIGNAL FA_lev5_col26_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col26_inst1_port_S: std_logic;
SIGNAL FA_lev5_col26_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col26_inst2_port_S: std_logic;
SIGNAL FA_lev5_col26_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col26_inst3_port_S: std_logic;
SIGNAL FA_lev5_col26_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col27_inst0_port_S: std_logic;
SIGNAL FA_lev5_col27_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col27_inst1_port_S: std_logic;
SIGNAL FA_lev5_col27_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col27_inst2_port_S: std_logic;
SIGNAL FA_lev5_col27_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col27_inst3_port_S: std_logic;
SIGNAL FA_lev5_col27_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col28_inst0_port_S: std_logic;
SIGNAL FA_lev5_col28_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col28_inst1_port_S: std_logic;
SIGNAL FA_lev5_col28_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col28_inst2_port_S: std_logic;
SIGNAL FA_lev5_col28_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col28_inst3_port_S: std_logic;
SIGNAL FA_lev5_col28_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col29_inst0_port_S: std_logic;
SIGNAL FA_lev5_col29_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col29_inst1_port_S: std_logic;
SIGNAL FA_lev5_col29_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col29_inst2_port_S: std_logic;
SIGNAL FA_lev5_col29_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col29_inst3_port_S: std_logic;
SIGNAL FA_lev5_col29_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col30_inst0_port_S: std_logic;
SIGNAL FA_lev5_col30_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col30_inst1_port_S: std_logic;
SIGNAL FA_lev5_col30_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col30_inst2_port_S: std_logic;
SIGNAL FA_lev5_col30_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col30_inst3_port_S: std_logic;
SIGNAL FA_lev5_col30_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col31_inst0_port_S: std_logic;
SIGNAL FA_lev5_col31_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col31_inst1_port_S: std_logic;
SIGNAL FA_lev5_col31_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col31_inst2_port_S: std_logic;
SIGNAL FA_lev5_col31_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col31_inst3_port_S: std_logic;
SIGNAL FA_lev5_col31_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col32_inst0_port_S: std_logic;
SIGNAL FA_lev5_col32_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col32_inst1_port_S: std_logic;
SIGNAL FA_lev5_col32_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col32_inst2_port_S: std_logic;
SIGNAL FA_lev5_col32_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col32_inst3_port_S: std_logic;
SIGNAL FA_lev5_col32_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col33_inst0_port_S: std_logic;
SIGNAL FA_lev5_col33_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col33_inst1_port_S: std_logic;
SIGNAL FA_lev5_col33_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col33_inst2_port_S: std_logic;
SIGNAL FA_lev5_col33_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col33_inst3_port_S: std_logic;
SIGNAL FA_lev5_col33_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col34_inst0_port_S: std_logic;
SIGNAL FA_lev5_col34_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col34_inst1_port_S: std_logic;
SIGNAL FA_lev5_col34_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col34_inst2_port_S: std_logic;
SIGNAL FA_lev5_col34_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col34_inst3_port_S: std_logic;
SIGNAL FA_lev5_col34_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col35_inst0_port_S: std_logic;
SIGNAL FA_lev5_col35_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col35_inst1_port_S: std_logic;
SIGNAL FA_lev5_col35_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col35_inst2_port_S: std_logic;
SIGNAL FA_lev5_col35_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col35_inst3_port_S: std_logic;
SIGNAL FA_lev5_col35_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col36_inst0_port_S: std_logic;
SIGNAL FA_lev5_col36_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col36_inst1_port_S: std_logic;
SIGNAL FA_lev5_col36_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col36_inst2_port_S: std_logic;
SIGNAL FA_lev5_col36_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col36_inst3_port_S: std_logic;
SIGNAL FA_lev5_col36_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col37_inst0_port_S: std_logic;
SIGNAL FA_lev5_col37_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col37_inst1_port_S: std_logic;
SIGNAL FA_lev5_col37_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col37_inst2_port_S: std_logic;
SIGNAL FA_lev5_col37_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col37_inst3_port_S: std_logic;
SIGNAL FA_lev5_col37_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col38_inst0_port_S: std_logic;
SIGNAL FA_lev5_col38_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col38_inst1_port_S: std_logic;
SIGNAL FA_lev5_col38_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col38_inst2_port_S: std_logic;
SIGNAL FA_lev5_col38_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col38_inst3_port_S: std_logic;
SIGNAL FA_lev5_col38_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col39_inst0_port_S: std_logic;
SIGNAL FA_lev5_col39_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col39_inst1_port_S: std_logic;
SIGNAL FA_lev5_col39_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col39_inst2_port_S: std_logic;
SIGNAL FA_lev5_col39_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col39_inst3_port_S: std_logic;
SIGNAL FA_lev5_col39_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col40_inst0_port_S: std_logic;
SIGNAL FA_lev5_col40_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col40_inst1_port_S: std_logic;
SIGNAL FA_lev5_col40_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col40_inst2_port_S: std_logic;
SIGNAL FA_lev5_col40_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col40_inst3_port_S: std_logic;
SIGNAL FA_lev5_col40_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col41_inst0_port_S: std_logic;
SIGNAL FA_lev5_col41_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col41_inst1_port_S: std_logic;
SIGNAL FA_lev5_col41_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col41_inst2_port_S: std_logic;
SIGNAL FA_lev5_col41_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col41_inst3_port_S: std_logic;
SIGNAL FA_lev5_col41_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col42_inst0_port_S: std_logic;
SIGNAL FA_lev5_col42_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col42_inst1_port_S: std_logic;
SIGNAL FA_lev5_col42_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col42_inst2_port_S: std_logic;
SIGNAL FA_lev5_col42_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col42_inst3_port_S: std_logic;
SIGNAL FA_lev5_col42_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col43_inst0_port_S: std_logic;
SIGNAL FA_lev5_col43_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col43_inst1_port_S: std_logic;
SIGNAL FA_lev5_col43_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col43_inst2_port_S: std_logic;
SIGNAL FA_lev5_col43_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col43_inst3_port_S: std_logic;
SIGNAL FA_lev5_col43_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col44_inst0_port_S: std_logic;
SIGNAL FA_lev5_col44_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col44_inst1_port_S: std_logic;
SIGNAL FA_lev5_col44_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col44_inst2_port_S: std_logic;
SIGNAL FA_lev5_col44_inst2_port_COUT: std_logic;
SIGNAL HA_lev5_col44_inst3_port_S: std_logic;
SIGNAL HA_lev5_col44_inst3_port_COUT: std_logic;
SIGNAL FA_lev5_col45_inst0_port_S: std_logic;
SIGNAL FA_lev5_col45_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col45_inst1_port_S: std_logic;
SIGNAL FA_lev5_col45_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col45_inst2_port_S: std_logic;
SIGNAL FA_lev5_col45_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col46_inst0_port_S: std_logic;
SIGNAL FA_lev5_col46_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col46_inst1_port_S: std_logic;
SIGNAL FA_lev5_col46_inst1_port_COUT: std_logic;
SIGNAL HA_lev5_col46_inst2_port_S: std_logic;
SIGNAL HA_lev5_col46_inst2_port_COUT: std_logic;
SIGNAL FA_lev5_col47_inst0_port_S: std_logic;
SIGNAL FA_lev5_col47_inst0_port_COUT: std_logic;
SIGNAL FA_lev5_col47_inst1_port_S: std_logic;
SIGNAL FA_lev5_col47_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col48_inst0_port_S: std_logic;
SIGNAL FA_lev5_col48_inst0_port_COUT: std_logic;
SIGNAL HA_lev5_col48_inst1_port_S: std_logic;
SIGNAL HA_lev5_col48_inst1_port_COUT: std_logic;
SIGNAL FA_lev5_col49_inst0_port_S: std_logic;
SIGNAL FA_lev5_col49_inst0_port_COUT: std_logic;
SIGNAL HA_lev5_col50_inst0_port_S: std_logic;
SIGNAL HA_lev5_col50_inst0_port_COUT: std_logic;
SIGNAL HA_lev4_col10_inst0_port_S: std_logic;
SIGNAL HA_lev4_col10_inst0_port_COUT: std_logic;
SIGNAL HA_lev4_col11_inst0_port_S: std_logic;
SIGNAL HA_lev4_col11_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col12_inst0_port_S: std_logic;
SIGNAL FA_lev4_col12_inst0_port_COUT: std_logic;
SIGNAL HA_lev4_col12_inst1_port_S: std_logic;
SIGNAL HA_lev4_col12_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col13_inst0_port_S: std_logic;
SIGNAL FA_lev4_col13_inst0_port_COUT: std_logic;
SIGNAL HA_lev4_col13_inst1_port_S: std_logic;
SIGNAL HA_lev4_col13_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col14_inst0_port_S: std_logic;
SIGNAL FA_lev4_col14_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col14_inst1_port_S: std_logic;
SIGNAL FA_lev4_col14_inst1_port_COUT: std_logic;
SIGNAL HA_lev4_col14_inst2_port_S: std_logic;
SIGNAL HA_lev4_col14_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col15_inst0_port_S: std_logic;
SIGNAL FA_lev4_col15_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col15_inst1_port_S: std_logic;
SIGNAL FA_lev4_col15_inst1_port_COUT: std_logic;
SIGNAL HA_lev4_col15_inst2_port_S: std_logic;
SIGNAL HA_lev4_col15_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col16_inst0_port_S: std_logic;
SIGNAL FA_lev4_col16_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col16_inst1_port_S: std_logic;
SIGNAL FA_lev4_col16_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col16_inst2_port_S: std_logic;
SIGNAL FA_lev4_col16_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col17_inst0_port_S: std_logic;
SIGNAL FA_lev4_col17_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col17_inst1_port_S: std_logic;
SIGNAL FA_lev4_col17_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col17_inst2_port_S: std_logic;
SIGNAL FA_lev4_col17_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col18_inst0_port_S: std_logic;
SIGNAL FA_lev4_col18_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col18_inst1_port_S: std_logic;
SIGNAL FA_lev4_col18_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col18_inst2_port_S: std_logic;
SIGNAL FA_lev4_col18_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col19_inst0_port_S: std_logic;
SIGNAL FA_lev4_col19_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col19_inst1_port_S: std_logic;
SIGNAL FA_lev4_col19_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col19_inst2_port_S: std_logic;
SIGNAL FA_lev4_col19_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col20_inst0_port_S: std_logic;
SIGNAL FA_lev4_col20_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col20_inst1_port_S: std_logic;
SIGNAL FA_lev4_col20_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col20_inst2_port_S: std_logic;
SIGNAL FA_lev4_col20_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col21_inst0_port_S: std_logic;
SIGNAL FA_lev4_col21_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col21_inst1_port_S: std_logic;
SIGNAL FA_lev4_col21_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col21_inst2_port_S: std_logic;
SIGNAL FA_lev4_col21_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col22_inst0_port_S: std_logic;
SIGNAL FA_lev4_col22_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col22_inst1_port_S: std_logic;
SIGNAL FA_lev4_col22_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col22_inst2_port_S: std_logic;
SIGNAL FA_lev4_col22_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col23_inst0_port_S: std_logic;
SIGNAL FA_lev4_col23_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col23_inst1_port_S: std_logic;
SIGNAL FA_lev4_col23_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col23_inst2_port_S: std_logic;
SIGNAL FA_lev4_col23_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col24_inst0_port_S: std_logic;
SIGNAL FA_lev4_col24_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col24_inst1_port_S: std_logic;
SIGNAL FA_lev4_col24_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col24_inst2_port_S: std_logic;
SIGNAL FA_lev4_col24_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col25_inst0_port_S: std_logic;
SIGNAL FA_lev4_col25_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col25_inst1_port_S: std_logic;
SIGNAL FA_lev4_col25_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col25_inst2_port_S: std_logic;
SIGNAL FA_lev4_col25_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col26_inst0_port_S: std_logic;
SIGNAL FA_lev4_col26_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col26_inst1_port_S: std_logic;
SIGNAL FA_lev4_col26_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col26_inst2_port_S: std_logic;
SIGNAL FA_lev4_col26_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col27_inst0_port_S: std_logic;
SIGNAL FA_lev4_col27_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col27_inst1_port_S: std_logic;
SIGNAL FA_lev4_col27_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col27_inst2_port_S: std_logic;
SIGNAL FA_lev4_col27_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col28_inst0_port_S: std_logic;
SIGNAL FA_lev4_col28_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col28_inst1_port_S: std_logic;
SIGNAL FA_lev4_col28_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col28_inst2_port_S: std_logic;
SIGNAL FA_lev4_col28_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col29_inst0_port_S: std_logic;
SIGNAL FA_lev4_col29_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col29_inst1_port_S: std_logic;
SIGNAL FA_lev4_col29_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col29_inst2_port_S: std_logic;
SIGNAL FA_lev4_col29_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col30_inst0_port_S: std_logic;
SIGNAL FA_lev4_col30_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col30_inst1_port_S: std_logic;
SIGNAL FA_lev4_col30_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col30_inst2_port_S: std_logic;
SIGNAL FA_lev4_col30_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col31_inst0_port_S: std_logic;
SIGNAL FA_lev4_col31_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col31_inst1_port_S: std_logic;
SIGNAL FA_lev4_col31_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col31_inst2_port_S: std_logic;
SIGNAL FA_lev4_col31_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col32_inst0_port_S: std_logic;
SIGNAL FA_lev4_col32_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col32_inst1_port_S: std_logic;
SIGNAL FA_lev4_col32_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col32_inst2_port_S: std_logic;
SIGNAL FA_lev4_col32_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col33_inst0_port_S: std_logic;
SIGNAL FA_lev4_col33_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col33_inst1_port_S: std_logic;
SIGNAL FA_lev4_col33_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col33_inst2_port_S: std_logic;
SIGNAL FA_lev4_col33_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col34_inst0_port_S: std_logic;
SIGNAL FA_lev4_col34_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col34_inst1_port_S: std_logic;
SIGNAL FA_lev4_col34_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col34_inst2_port_S: std_logic;
SIGNAL FA_lev4_col34_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col35_inst0_port_S: std_logic;
SIGNAL FA_lev4_col35_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col35_inst1_port_S: std_logic;
SIGNAL FA_lev4_col35_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col35_inst2_port_S: std_logic;
SIGNAL FA_lev4_col35_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col36_inst0_port_S: std_logic;
SIGNAL FA_lev4_col36_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col36_inst1_port_S: std_logic;
SIGNAL FA_lev4_col36_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col36_inst2_port_S: std_logic;
SIGNAL FA_lev4_col36_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col37_inst0_port_S: std_logic;
SIGNAL FA_lev4_col37_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col37_inst1_port_S: std_logic;
SIGNAL FA_lev4_col37_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col37_inst2_port_S: std_logic;
SIGNAL FA_lev4_col37_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col38_inst0_port_S: std_logic;
SIGNAL FA_lev4_col38_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col38_inst1_port_S: std_logic;
SIGNAL FA_lev4_col38_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col38_inst2_port_S: std_logic;
SIGNAL FA_lev4_col38_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col39_inst0_port_S: std_logic;
SIGNAL FA_lev4_col39_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col39_inst1_port_S: std_logic;
SIGNAL FA_lev4_col39_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col39_inst2_port_S: std_logic;
SIGNAL FA_lev4_col39_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col40_inst0_port_S: std_logic;
SIGNAL FA_lev4_col40_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col40_inst1_port_S: std_logic;
SIGNAL FA_lev4_col40_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col40_inst2_port_S: std_logic;
SIGNAL FA_lev4_col40_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col41_inst0_port_S: std_logic;
SIGNAL FA_lev4_col41_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col41_inst1_port_S: std_logic;
SIGNAL FA_lev4_col41_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col41_inst2_port_S: std_logic;
SIGNAL FA_lev4_col41_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col42_inst0_port_S: std_logic;
SIGNAL FA_lev4_col42_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col42_inst1_port_S: std_logic;
SIGNAL FA_lev4_col42_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col42_inst2_port_S: std_logic;
SIGNAL FA_lev4_col42_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col43_inst0_port_S: std_logic;
SIGNAL FA_lev4_col43_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col43_inst1_port_S: std_logic;
SIGNAL FA_lev4_col43_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col43_inst2_port_S: std_logic;
SIGNAL FA_lev4_col43_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col44_inst0_port_S: std_logic;
SIGNAL FA_lev4_col44_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col44_inst1_port_S: std_logic;
SIGNAL FA_lev4_col44_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col44_inst2_port_S: std_logic;
SIGNAL FA_lev4_col44_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col45_inst0_port_S: std_logic;
SIGNAL FA_lev4_col45_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col45_inst1_port_S: std_logic;
SIGNAL FA_lev4_col45_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col45_inst2_port_S: std_logic;
SIGNAL FA_lev4_col45_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col46_inst0_port_S: std_logic;
SIGNAL FA_lev4_col46_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col46_inst1_port_S: std_logic;
SIGNAL FA_lev4_col46_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col46_inst2_port_S: std_logic;
SIGNAL FA_lev4_col46_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col47_inst0_port_S: std_logic;
SIGNAL FA_lev4_col47_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col47_inst1_port_S: std_logic;
SIGNAL FA_lev4_col47_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col47_inst2_port_S: std_logic;
SIGNAL FA_lev4_col47_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col48_inst0_port_S: std_logic;
SIGNAL FA_lev4_col48_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col48_inst1_port_S: std_logic;
SIGNAL FA_lev4_col48_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col48_inst2_port_S: std_logic;
SIGNAL FA_lev4_col48_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col49_inst0_port_S: std_logic;
SIGNAL FA_lev4_col49_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col49_inst1_port_S: std_logic;
SIGNAL FA_lev4_col49_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col49_inst2_port_S: std_logic;
SIGNAL FA_lev4_col49_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col50_inst0_port_S: std_logic;
SIGNAL FA_lev4_col50_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col50_inst1_port_S: std_logic;
SIGNAL FA_lev4_col50_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col50_inst2_port_S: std_logic;
SIGNAL FA_lev4_col50_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col51_inst0_port_S: std_logic;
SIGNAL FA_lev4_col51_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col51_inst1_port_S: std_logic;
SIGNAL FA_lev4_col51_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col51_inst2_port_S: std_logic;
SIGNAL FA_lev4_col51_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col52_inst0_port_S: std_logic;
SIGNAL FA_lev4_col52_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col52_inst1_port_S: std_logic;
SIGNAL FA_lev4_col52_inst1_port_COUT: std_logic;
SIGNAL HA_lev4_col52_inst2_port_S: std_logic;
SIGNAL HA_lev4_col52_inst2_port_COUT: std_logic;
SIGNAL FA_lev4_col53_inst0_port_S: std_logic;
SIGNAL FA_lev4_col53_inst0_port_COUT: std_logic;
SIGNAL FA_lev4_col53_inst1_port_S: std_logic;
SIGNAL FA_lev4_col53_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col54_inst0_port_S: std_logic;
SIGNAL FA_lev4_col54_inst0_port_COUT: std_logic;
SIGNAL HA_lev4_col54_inst1_port_S: std_logic;
SIGNAL HA_lev4_col54_inst1_port_COUT: std_logic;
SIGNAL FA_lev4_col55_inst0_port_S: std_logic;
SIGNAL FA_lev4_col55_inst0_port_COUT: std_logic;
SIGNAL HA_lev4_col56_inst0_port_S: std_logic;
SIGNAL HA_lev4_col56_inst0_port_COUT: std_logic;
SIGNAL HA_lev3_col6_inst0_port_S: std_logic;
SIGNAL HA_lev3_col6_inst0_port_COUT: std_logic;
SIGNAL HA_lev3_col7_inst0_port_S: std_logic;
SIGNAL HA_lev3_col7_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col8_inst0_port_S: std_logic;
SIGNAL FA_lev3_col8_inst0_port_COUT: std_logic;
SIGNAL HA_lev3_col8_inst1_port_S: std_logic;
SIGNAL HA_lev3_col8_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col9_inst0_port_S: std_logic;
SIGNAL FA_lev3_col9_inst0_port_COUT: std_logic;
SIGNAL HA_lev3_col9_inst1_port_S: std_logic;
SIGNAL HA_lev3_col9_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col10_inst0_port_S: std_logic;
SIGNAL FA_lev3_col10_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col10_inst1_port_S: std_logic;
SIGNAL FA_lev3_col10_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col11_inst0_port_S: std_logic;
SIGNAL FA_lev3_col11_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col11_inst1_port_S: std_logic;
SIGNAL FA_lev3_col11_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col12_inst0_port_S: std_logic;
SIGNAL FA_lev3_col12_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col12_inst1_port_S: std_logic;
SIGNAL FA_lev3_col12_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col13_inst0_port_S: std_logic;
SIGNAL FA_lev3_col13_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col13_inst1_port_S: std_logic;
SIGNAL FA_lev3_col13_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col14_inst0_port_S: std_logic;
SIGNAL FA_lev3_col14_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col14_inst1_port_S: std_logic;
SIGNAL FA_lev3_col14_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col15_inst0_port_S: std_logic;
SIGNAL FA_lev3_col15_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col15_inst1_port_S: std_logic;
SIGNAL FA_lev3_col15_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col16_inst0_port_S: std_logic;
SIGNAL FA_lev3_col16_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col16_inst1_port_S: std_logic;
SIGNAL FA_lev3_col16_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col17_inst0_port_S: std_logic;
SIGNAL FA_lev3_col17_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col17_inst1_port_S: std_logic;
SIGNAL FA_lev3_col17_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col18_inst0_port_S: std_logic;
SIGNAL FA_lev3_col18_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col18_inst1_port_S: std_logic;
SIGNAL FA_lev3_col18_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col19_inst0_port_S: std_logic;
SIGNAL FA_lev3_col19_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col19_inst1_port_S: std_logic;
SIGNAL FA_lev3_col19_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col20_inst0_port_S: std_logic;
SIGNAL FA_lev3_col20_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col20_inst1_port_S: std_logic;
SIGNAL FA_lev3_col20_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col21_inst0_port_S: std_logic;
SIGNAL FA_lev3_col21_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col21_inst1_port_S: std_logic;
SIGNAL FA_lev3_col21_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col22_inst0_port_S: std_logic;
SIGNAL FA_lev3_col22_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col22_inst1_port_S: std_logic;
SIGNAL FA_lev3_col22_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col23_inst0_port_S: std_logic;
SIGNAL FA_lev3_col23_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col23_inst1_port_S: std_logic;
SIGNAL FA_lev3_col23_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col24_inst0_port_S: std_logic;
SIGNAL FA_lev3_col24_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col24_inst1_port_S: std_logic;
SIGNAL FA_lev3_col24_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col25_inst0_port_S: std_logic;
SIGNAL FA_lev3_col25_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col25_inst1_port_S: std_logic;
SIGNAL FA_lev3_col25_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col26_inst0_port_S: std_logic;
SIGNAL FA_lev3_col26_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col26_inst1_port_S: std_logic;
SIGNAL FA_lev3_col26_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col27_inst0_port_S: std_logic;
SIGNAL FA_lev3_col27_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col27_inst1_port_S: std_logic;
SIGNAL FA_lev3_col27_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col28_inst0_port_S: std_logic;
SIGNAL FA_lev3_col28_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col28_inst1_port_S: std_logic;
SIGNAL FA_lev3_col28_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col29_inst0_port_S: std_logic;
SIGNAL FA_lev3_col29_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col29_inst1_port_S: std_logic;
SIGNAL FA_lev3_col29_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col30_inst0_port_S: std_logic;
SIGNAL FA_lev3_col30_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col30_inst1_port_S: std_logic;
SIGNAL FA_lev3_col30_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col31_inst0_port_S: std_logic;
SIGNAL FA_lev3_col31_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col31_inst1_port_S: std_logic;
SIGNAL FA_lev3_col31_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col32_inst0_port_S: std_logic;
SIGNAL FA_lev3_col32_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col32_inst1_port_S: std_logic;
SIGNAL FA_lev3_col32_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col33_inst0_port_S: std_logic;
SIGNAL FA_lev3_col33_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col33_inst1_port_S: std_logic;
SIGNAL FA_lev3_col33_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col34_inst0_port_S: std_logic;
SIGNAL FA_lev3_col34_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col34_inst1_port_S: std_logic;
SIGNAL FA_lev3_col34_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col35_inst0_port_S: std_logic;
SIGNAL FA_lev3_col35_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col35_inst1_port_S: std_logic;
SIGNAL FA_lev3_col35_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col36_inst0_port_S: std_logic;
SIGNAL FA_lev3_col36_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col36_inst1_port_S: std_logic;
SIGNAL FA_lev3_col36_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col37_inst0_port_S: std_logic;
SIGNAL FA_lev3_col37_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col37_inst1_port_S: std_logic;
SIGNAL FA_lev3_col37_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col38_inst0_port_S: std_logic;
SIGNAL FA_lev3_col38_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col38_inst1_port_S: std_logic;
SIGNAL FA_lev3_col38_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col39_inst0_port_S: std_logic;
SIGNAL FA_lev3_col39_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col39_inst1_port_S: std_logic;
SIGNAL FA_lev3_col39_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col40_inst0_port_S: std_logic;
SIGNAL FA_lev3_col40_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col40_inst1_port_S: std_logic;
SIGNAL FA_lev3_col40_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col41_inst0_port_S: std_logic;
SIGNAL FA_lev3_col41_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col41_inst1_port_S: std_logic;
SIGNAL FA_lev3_col41_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col42_inst0_port_S: std_logic;
SIGNAL FA_lev3_col42_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col42_inst1_port_S: std_logic;
SIGNAL FA_lev3_col42_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col43_inst0_port_S: std_logic;
SIGNAL FA_lev3_col43_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col43_inst1_port_S: std_logic;
SIGNAL FA_lev3_col43_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col44_inst0_port_S: std_logic;
SIGNAL FA_lev3_col44_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col44_inst1_port_S: std_logic;
SIGNAL FA_lev3_col44_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col45_inst0_port_S: std_logic;
SIGNAL FA_lev3_col45_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col45_inst1_port_S: std_logic;
SIGNAL FA_lev3_col45_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col46_inst0_port_S: std_logic;
SIGNAL FA_lev3_col46_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col46_inst1_port_S: std_logic;
SIGNAL FA_lev3_col46_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col47_inst0_port_S: std_logic;
SIGNAL FA_lev3_col47_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col47_inst1_port_S: std_logic;
SIGNAL FA_lev3_col47_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col48_inst0_port_S: std_logic;
SIGNAL FA_lev3_col48_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col48_inst1_port_S: std_logic;
SIGNAL FA_lev3_col48_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col49_inst0_port_S: std_logic;
SIGNAL FA_lev3_col49_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col49_inst1_port_S: std_logic;
SIGNAL FA_lev3_col49_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col50_inst0_port_S: std_logic;
SIGNAL FA_lev3_col50_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col50_inst1_port_S: std_logic;
SIGNAL FA_lev3_col50_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col51_inst0_port_S: std_logic;
SIGNAL FA_lev3_col51_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col51_inst1_port_S: std_logic;
SIGNAL FA_lev3_col51_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col52_inst0_port_S: std_logic;
SIGNAL FA_lev3_col52_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col52_inst1_port_S: std_logic;
SIGNAL FA_lev3_col52_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col53_inst0_port_S: std_logic;
SIGNAL FA_lev3_col53_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col53_inst1_port_S: std_logic;
SIGNAL FA_lev3_col53_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col54_inst0_port_S: std_logic;
SIGNAL FA_lev3_col54_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col54_inst1_port_S: std_logic;
SIGNAL FA_lev3_col54_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col55_inst0_port_S: std_logic;
SIGNAL FA_lev3_col55_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col55_inst1_port_S: std_logic;
SIGNAL FA_lev3_col55_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col56_inst0_port_S: std_logic;
SIGNAL FA_lev3_col56_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col56_inst1_port_S: std_logic;
SIGNAL FA_lev3_col56_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col57_inst0_port_S: std_logic;
SIGNAL FA_lev3_col57_inst0_port_COUT: std_logic;
SIGNAL FA_lev3_col57_inst1_port_S: std_logic;
SIGNAL FA_lev3_col57_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col58_inst0_port_S: std_logic;
SIGNAL FA_lev3_col58_inst0_port_COUT: std_logic;
SIGNAL HA_lev3_col58_inst1_port_S: std_logic;
SIGNAL HA_lev3_col58_inst1_port_COUT: std_logic;
SIGNAL FA_lev3_col59_inst0_port_S: std_logic;
SIGNAL FA_lev3_col59_inst0_port_COUT: std_logic;
SIGNAL HA_lev3_col60_inst0_port_S: std_logic;
SIGNAL HA_lev3_col60_inst0_port_COUT: std_logic;
SIGNAL HA_lev2_col4_inst0_port_S: std_logic;
SIGNAL HA_lev2_col4_inst0_port_COUT: std_logic;
SIGNAL HA_lev2_col5_inst0_port_S: std_logic;
SIGNAL HA_lev2_col5_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col6_inst0_port_S: std_logic;
SIGNAL FA_lev2_col6_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col7_inst0_port_S: std_logic;
SIGNAL FA_lev2_col7_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col8_inst0_port_S: std_logic;
SIGNAL FA_lev2_col8_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col9_inst0_port_S: std_logic;
SIGNAL FA_lev2_col9_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col10_inst0_port_S: std_logic;
SIGNAL FA_lev2_col10_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col11_inst0_port_S: std_logic;
SIGNAL FA_lev2_col11_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col12_inst0_port_S: std_logic;
SIGNAL FA_lev2_col12_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col13_inst0_port_S: std_logic;
SIGNAL FA_lev2_col13_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col14_inst0_port_S: std_logic;
SIGNAL FA_lev2_col14_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col15_inst0_port_S: std_logic;
SIGNAL FA_lev2_col15_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col16_inst0_port_S: std_logic;
SIGNAL FA_lev2_col16_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col17_inst0_port_S: std_logic;
SIGNAL FA_lev2_col17_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col18_inst0_port_S: std_logic;
SIGNAL FA_lev2_col18_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col19_inst0_port_S: std_logic;
SIGNAL FA_lev2_col19_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col20_inst0_port_S: std_logic;
SIGNAL FA_lev2_col20_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col21_inst0_port_S: std_logic;
SIGNAL FA_lev2_col21_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col22_inst0_port_S: std_logic;
SIGNAL FA_lev2_col22_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col23_inst0_port_S: std_logic;
SIGNAL FA_lev2_col23_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col24_inst0_port_S: std_logic;
SIGNAL FA_lev2_col24_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col25_inst0_port_S: std_logic;
SIGNAL FA_lev2_col25_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col26_inst0_port_S: std_logic;
SIGNAL FA_lev2_col26_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col27_inst0_port_S: std_logic;
SIGNAL FA_lev2_col27_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col28_inst0_port_S: std_logic;
SIGNAL FA_lev2_col28_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col29_inst0_port_S: std_logic;
SIGNAL FA_lev2_col29_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col30_inst0_port_S: std_logic;
SIGNAL FA_lev2_col30_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col31_inst0_port_S: std_logic;
SIGNAL FA_lev2_col31_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col32_inst0_port_S: std_logic;
SIGNAL FA_lev2_col32_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col33_inst0_port_S: std_logic;
SIGNAL FA_lev2_col33_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col34_inst0_port_S: std_logic;
SIGNAL FA_lev2_col34_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col35_inst0_port_S: std_logic;
SIGNAL FA_lev2_col35_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col36_inst0_port_S: std_logic;
SIGNAL FA_lev2_col36_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col37_inst0_port_S: std_logic;
SIGNAL FA_lev2_col37_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col38_inst0_port_S: std_logic;
SIGNAL FA_lev2_col38_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col39_inst0_port_S: std_logic;
SIGNAL FA_lev2_col39_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col40_inst0_port_S: std_logic;
SIGNAL FA_lev2_col40_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col41_inst0_port_S: std_logic;
SIGNAL FA_lev2_col41_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col42_inst0_port_S: std_logic;
SIGNAL FA_lev2_col42_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col43_inst0_port_S: std_logic;
SIGNAL FA_lev2_col43_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col44_inst0_port_S: std_logic;
SIGNAL FA_lev2_col44_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col45_inst0_port_S: std_logic;
SIGNAL FA_lev2_col45_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col46_inst0_port_S: std_logic;
SIGNAL FA_lev2_col46_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col47_inst0_port_S: std_logic;
SIGNAL FA_lev2_col47_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col48_inst0_port_S: std_logic;
SIGNAL FA_lev2_col48_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col49_inst0_port_S: std_logic;
SIGNAL FA_lev2_col49_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col50_inst0_port_S: std_logic;
SIGNAL FA_lev2_col50_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col51_inst0_port_S: std_logic;
SIGNAL FA_lev2_col51_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col52_inst0_port_S: std_logic;
SIGNAL FA_lev2_col52_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col53_inst0_port_S: std_logic;
SIGNAL FA_lev2_col53_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col54_inst0_port_S: std_logic;
SIGNAL FA_lev2_col54_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col55_inst0_port_S: std_logic;
SIGNAL FA_lev2_col55_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col56_inst0_port_S: std_logic;
SIGNAL FA_lev2_col56_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col57_inst0_port_S: std_logic;
SIGNAL FA_lev2_col57_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col58_inst0_port_S: std_logic;
SIGNAL FA_lev2_col58_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col59_inst0_port_S: std_logic;
SIGNAL FA_lev2_col59_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col60_inst0_port_S: std_logic;
SIGNAL FA_lev2_col60_inst0_port_COUT: std_logic;
SIGNAL FA_lev2_col61_inst0_port_S: std_logic;
SIGNAL FA_lev2_col61_inst0_port_COUT: std_logic;
SIGNAL HA_lev2_col62_inst0_port_S: std_logic;
SIGNAL HA_lev2_col62_inst0_port_COUT: std_logic;
SIGNAL HA_lev1_col2_inst0_port_S: std_logic;
SIGNAL HA_lev1_col2_inst0_port_COUT: std_logic;
SIGNAL HA_lev1_col3_inst0_port_S: std_logic;
SIGNAL HA_lev1_col3_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col4_inst0_port_S: std_logic;
SIGNAL FA_lev1_col4_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col5_inst0_port_S: std_logic;
SIGNAL FA_lev1_col5_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col6_inst0_port_S: std_logic;
SIGNAL FA_lev1_col6_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col7_inst0_port_S: std_logic;
SIGNAL FA_lev1_col7_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col8_inst0_port_S: std_logic;
SIGNAL FA_lev1_col8_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col9_inst0_port_S: std_logic;
SIGNAL FA_lev1_col9_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col10_inst0_port_S: std_logic;
SIGNAL FA_lev1_col10_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col11_inst0_port_S: std_logic;
SIGNAL FA_lev1_col11_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col12_inst0_port_S: std_logic;
SIGNAL FA_lev1_col12_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col13_inst0_port_S: std_logic;
SIGNAL FA_lev1_col13_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col14_inst0_port_S: std_logic;
SIGNAL FA_lev1_col14_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col15_inst0_port_S: std_logic;
SIGNAL FA_lev1_col15_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col16_inst0_port_S: std_logic;
SIGNAL FA_lev1_col16_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col17_inst0_port_S: std_logic;
SIGNAL FA_lev1_col17_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col18_inst0_port_S: std_logic;
SIGNAL FA_lev1_col18_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col19_inst0_port_S: std_logic;
SIGNAL FA_lev1_col19_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col20_inst0_port_S: std_logic;
SIGNAL FA_lev1_col20_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col21_inst0_port_S: std_logic;
SIGNAL FA_lev1_col21_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col22_inst0_port_S: std_logic;
SIGNAL FA_lev1_col22_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col23_inst0_port_S: std_logic;
SIGNAL FA_lev1_col23_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col24_inst0_port_S: std_logic;
SIGNAL FA_lev1_col24_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col25_inst0_port_S: std_logic;
SIGNAL FA_lev1_col25_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col26_inst0_port_S: std_logic;
SIGNAL FA_lev1_col26_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col27_inst0_port_S: std_logic;
SIGNAL FA_lev1_col27_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col28_inst0_port_S: std_logic;
SIGNAL FA_lev1_col28_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col29_inst0_port_S: std_logic;
SIGNAL FA_lev1_col29_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col30_inst0_port_S: std_logic;
SIGNAL FA_lev1_col30_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col31_inst0_port_S: std_logic;
SIGNAL FA_lev1_col31_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col32_inst0_port_S: std_logic;
SIGNAL FA_lev1_col32_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col33_inst0_port_S: std_logic;
SIGNAL FA_lev1_col33_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col34_inst0_port_S: std_logic;
SIGNAL FA_lev1_col34_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col35_inst0_port_S: std_logic;
SIGNAL FA_lev1_col35_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col36_inst0_port_S: std_logic;
SIGNAL FA_lev1_col36_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col37_inst0_port_S: std_logic;
SIGNAL FA_lev1_col37_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col38_inst0_port_S: std_logic;
SIGNAL FA_lev1_col38_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col39_inst0_port_S: std_logic;
SIGNAL FA_lev1_col39_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col40_inst0_port_S: std_logic;
SIGNAL FA_lev1_col40_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col41_inst0_port_S: std_logic;
SIGNAL FA_lev1_col41_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col42_inst0_port_S: std_logic;
SIGNAL FA_lev1_col42_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col43_inst0_port_S: std_logic;
SIGNAL FA_lev1_col43_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col44_inst0_port_S: std_logic;
SIGNAL FA_lev1_col44_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col45_inst0_port_S: std_logic;
SIGNAL FA_lev1_col45_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col46_inst0_port_S: std_logic;
SIGNAL FA_lev1_col46_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col47_inst0_port_S: std_logic;
SIGNAL FA_lev1_col47_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col48_inst0_port_S: std_logic;
SIGNAL FA_lev1_col48_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col49_inst0_port_S: std_logic;
SIGNAL FA_lev1_col49_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col50_inst0_port_S: std_logic;
SIGNAL FA_lev1_col50_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col51_inst0_port_S: std_logic;
SIGNAL FA_lev1_col51_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col52_inst0_port_S: std_logic;
SIGNAL FA_lev1_col52_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col53_inst0_port_S: std_logic;
SIGNAL FA_lev1_col53_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col54_inst0_port_S: std_logic;
SIGNAL FA_lev1_col54_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col55_inst0_port_S: std_logic;
SIGNAL FA_lev1_col55_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col56_inst0_port_S: std_logic;
SIGNAL FA_lev1_col56_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col57_inst0_port_S: std_logic;
SIGNAL FA_lev1_col57_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col58_inst0_port_S: std_logic;
SIGNAL FA_lev1_col58_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col59_inst0_port_S: std_logic;
SIGNAL FA_lev1_col59_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col60_inst0_port_S: std_logic;
SIGNAL FA_lev1_col60_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col61_inst0_port_S: std_logic;
SIGNAL FA_lev1_col61_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col62_inst0_port_S: std_logic;
SIGNAL FA_lev1_col62_inst0_port_COUT: std_logic;
SIGNAL FA_lev1_col63_inst0_port_S: std_logic;
SIGNAL FA_lev1_col63_inst0_port_COUT: std_logic;

BEGIN

-- Level no 7
HA_lev6_col24_inst0: HA PORT MAP(PP_IN(0)(24), PP_IN(1)(24), HA_lev6_col24_inst0_port_S, HA_lev6_col24_inst0_port_COUT);
HA_lev6_col25_inst0: HA PORT MAP(PP_IN(0)(25), PP_IN(1)(25), HA_lev6_col25_inst0_port_S, HA_lev6_col25_inst0_port_COUT);
FA_lev6_col26_inst0: FA PORT MAP(PP_IN(0)(26), PP_IN(1)(26), PP_IN(2)(26), FA_lev6_col26_inst0_port_S, FA_lev6_col26_inst0_port_COUT);
HA_lev6_col26_inst1: HA PORT MAP(PP_IN(3)(26), PP_IN(4)(26), HA_lev6_col26_inst1_port_S, HA_lev6_col26_inst1_port_COUT);
FA_lev6_col27_inst0: FA PORT MAP(PP_IN(0)(27), PP_IN(1)(27), PP_IN(2)(27), FA_lev6_col27_inst0_port_S, FA_lev6_col27_inst0_port_COUT);
HA_lev6_col27_inst1: HA PORT MAP(PP_IN(3)(27), PP_IN(4)(27), HA_lev6_col27_inst1_port_S, HA_lev6_col27_inst1_port_COUT);
FA_lev6_col28_inst0: FA PORT MAP(PP_IN(0)(28), PP_IN(1)(28), PP_IN(2)(28), FA_lev6_col28_inst0_port_S, FA_lev6_col28_inst0_port_COUT);
FA_lev6_col28_inst1: FA PORT MAP(PP_IN(3)(28), PP_IN(4)(28), PP_IN(5)(28), FA_lev6_col28_inst1_port_S, FA_lev6_col28_inst1_port_COUT);
HA_lev6_col28_inst2: HA PORT MAP(PP_IN(6)(28), PP_IN(7)(28), HA_lev6_col28_inst2_port_S, HA_lev6_col28_inst2_port_COUT);
FA_lev6_col29_inst0: FA PORT MAP(PP_IN(0)(29), PP_IN(1)(29), PP_IN(2)(29), FA_lev6_col29_inst0_port_S, FA_lev6_col29_inst0_port_COUT);
FA_lev6_col29_inst1: FA PORT MAP(PP_IN(3)(29), PP_IN(4)(29), PP_IN(5)(29), FA_lev6_col29_inst1_port_S, FA_lev6_col29_inst1_port_COUT);
HA_lev6_col29_inst2: HA PORT MAP(PP_IN(6)(29), PP_IN(7)(29), HA_lev6_col29_inst2_port_S, HA_lev6_col29_inst2_port_COUT);
FA_lev6_col30_inst0: FA PORT MAP(PP_IN(0)(30), PP_IN(1)(30), PP_IN(2)(30), FA_lev6_col30_inst0_port_S, FA_lev6_col30_inst0_port_COUT);
FA_lev6_col30_inst1: FA PORT MAP(PP_IN(3)(30), PP_IN(4)(30), PP_IN(5)(30), FA_lev6_col30_inst1_port_S, FA_lev6_col30_inst1_port_COUT);
FA_lev6_col30_inst2: FA PORT MAP(PP_IN(6)(30), PP_IN(7)(30), PP_IN(8)(30), FA_lev6_col30_inst2_port_S, FA_lev6_col30_inst2_port_COUT);
HA_lev6_col30_inst3: HA PORT MAP(PP_IN(9)(30), PP_IN(10)(30), HA_lev6_col30_inst3_port_S, HA_lev6_col30_inst3_port_COUT);
FA_lev6_col31_inst0: FA PORT MAP(PP_IN(0)(31), PP_IN(1)(31), PP_IN(2)(31), FA_lev6_col31_inst0_port_S, FA_lev6_col31_inst0_port_COUT);
FA_lev6_col31_inst1: FA PORT MAP(PP_IN(3)(31), PP_IN(4)(31), PP_IN(5)(31), FA_lev6_col31_inst1_port_S, FA_lev6_col31_inst1_port_COUT);
FA_lev6_col31_inst2: FA PORT MAP(PP_IN(6)(31), PP_IN(7)(31), PP_IN(8)(31), FA_lev6_col31_inst2_port_S, FA_lev6_col31_inst2_port_COUT);
HA_lev6_col31_inst3: HA PORT MAP(PP_IN(9)(31), PP_IN(10)(31), HA_lev6_col31_inst3_port_S, HA_lev6_col31_inst3_port_COUT);
FA_lev6_col32_inst0: FA PORT MAP(PP_IN(0)(32), PP_IN(1)(32), PP_IN(2)(32), FA_lev6_col32_inst0_port_S, FA_lev6_col32_inst0_port_COUT);
FA_lev6_col32_inst1: FA PORT MAP(PP_IN(3)(32), PP_IN(4)(32), PP_IN(5)(32), FA_lev6_col32_inst1_port_S, FA_lev6_col32_inst1_port_COUT);
FA_lev6_col32_inst2: FA PORT MAP(PP_IN(6)(32), PP_IN(7)(32), PP_IN(8)(32), FA_lev6_col32_inst2_port_S, FA_lev6_col32_inst2_port_COUT);
FA_lev6_col32_inst3: FA PORT MAP(PP_IN(9)(32), PP_IN(10)(32), PP_IN(11)(32), FA_lev6_col32_inst3_port_S, FA_lev6_col32_inst3_port_COUT);
FA_lev6_col33_inst0: FA PORT MAP(PP_IN(0)(33), PP_IN(1)(33), PP_IN(2)(33), FA_lev6_col33_inst0_port_S, FA_lev6_col33_inst0_port_COUT);
FA_lev6_col33_inst1: FA PORT MAP(PP_IN(3)(33), PP_IN(4)(33), PP_IN(5)(33), FA_lev6_col33_inst1_port_S, FA_lev6_col33_inst1_port_COUT);
FA_lev6_col33_inst2: FA PORT MAP(PP_IN(6)(33), PP_IN(7)(33), PP_IN(8)(33), FA_lev6_col33_inst2_port_S, FA_lev6_col33_inst2_port_COUT);
FA_lev6_col33_inst3: FA PORT MAP(PP_IN(9)(33), PP_IN(10)(33), PP_IN(11)(33), FA_lev6_col33_inst3_port_S, FA_lev6_col33_inst3_port_COUT);
FA_lev6_col34_inst0: FA PORT MAP(PP_IN(0)(34), PP_IN(1)(34), PP_IN(2)(34), FA_lev6_col34_inst0_port_S, FA_lev6_col34_inst0_port_COUT);
FA_lev6_col34_inst1: FA PORT MAP(PP_IN(3)(34), PP_IN(4)(34), PP_IN(5)(34), FA_lev6_col34_inst1_port_S, FA_lev6_col34_inst1_port_COUT);
FA_lev6_col34_inst2: FA PORT MAP(PP_IN(6)(34), PP_IN(7)(34), PP_IN(8)(34), FA_lev6_col34_inst2_port_S, FA_lev6_col34_inst2_port_COUT);
FA_lev6_col34_inst3: FA PORT MAP(PP_IN(9)(34), PP_IN(10)(34), PP_IN(11)(34), FA_lev6_col34_inst3_port_S, FA_lev6_col34_inst3_port_COUT);
FA_lev6_col35_inst0: FA PORT MAP(PP_IN(0)(35), PP_IN(1)(35), PP_IN(2)(35), FA_lev6_col35_inst0_port_S, FA_lev6_col35_inst0_port_COUT);
FA_lev6_col35_inst1: FA PORT MAP(PP_IN(3)(35), PP_IN(4)(35), PP_IN(5)(35), FA_lev6_col35_inst1_port_S, FA_lev6_col35_inst1_port_COUT);
FA_lev6_col35_inst2: FA PORT MAP(PP_IN(6)(35), PP_IN(7)(35), PP_IN(8)(35), FA_lev6_col35_inst2_port_S, FA_lev6_col35_inst2_port_COUT);
FA_lev6_col35_inst3: FA PORT MAP(PP_IN(9)(35), PP_IN(10)(35), PP_IN(11)(35), FA_lev6_col35_inst3_port_S, FA_lev6_col35_inst3_port_COUT);
FA_lev6_col36_inst0: FA PORT MAP(PP_IN(0)(36), PP_IN(1)(36), PP_IN(2)(36), FA_lev6_col36_inst0_port_S, FA_lev6_col36_inst0_port_COUT);
FA_lev6_col36_inst1: FA PORT MAP(PP_IN(3)(36), PP_IN(4)(36), PP_IN(5)(36), FA_lev6_col36_inst1_port_S, FA_lev6_col36_inst1_port_COUT);
FA_lev6_col36_inst2: FA PORT MAP(PP_IN(6)(36), PP_IN(7)(36), PP_IN(8)(36), FA_lev6_col36_inst2_port_S, FA_lev6_col36_inst2_port_COUT);
HA_lev6_col36_inst3: HA PORT MAP(PP_IN(9)(36), PP_IN(10)(36), HA_lev6_col36_inst3_port_S, HA_lev6_col36_inst3_port_COUT);
FA_lev6_col37_inst0: FA PORT MAP(PP_IN(0)(37), PP_IN(1)(37), PP_IN(2)(37), FA_lev6_col37_inst0_port_S, FA_lev6_col37_inst0_port_COUT);
FA_lev6_col37_inst1: FA PORT MAP(PP_IN(3)(37), PP_IN(4)(37), PP_IN(5)(37), FA_lev6_col37_inst1_port_S, FA_lev6_col37_inst1_port_COUT);
FA_lev6_col37_inst2: FA PORT MAP(PP_IN(6)(37), PP_IN(7)(37), PP_IN(8)(37), FA_lev6_col37_inst2_port_S, FA_lev6_col37_inst2_port_COUT);
FA_lev6_col38_inst0: FA PORT MAP(PP_IN(0)(38), PP_IN(1)(38), PP_IN(2)(38), FA_lev6_col38_inst0_port_S, FA_lev6_col38_inst0_port_COUT);
FA_lev6_col38_inst1: FA PORT MAP(PP_IN(3)(38), PP_IN(4)(38), PP_IN(5)(38), FA_lev6_col38_inst1_port_S, FA_lev6_col38_inst1_port_COUT);
HA_lev6_col38_inst2: HA PORT MAP(PP_IN(6)(38), PP_IN(7)(38), HA_lev6_col38_inst2_port_S, HA_lev6_col38_inst2_port_COUT);
FA_lev6_col39_inst0: FA PORT MAP(PP_IN(0)(39), PP_IN(1)(39), PP_IN(2)(39), FA_lev6_col39_inst0_port_S, FA_lev6_col39_inst0_port_COUT);
FA_lev6_col39_inst1: FA PORT MAP(PP_IN(3)(39), PP_IN(4)(39), PP_IN(5)(39), FA_lev6_col39_inst1_port_S, FA_lev6_col39_inst1_port_COUT);
FA_lev6_col40_inst0: FA PORT MAP(PP_IN(0)(40), PP_IN(1)(40), PP_IN(2)(40), FA_lev6_col40_inst0_port_S, FA_lev6_col40_inst0_port_COUT);
HA_lev6_col40_inst1: HA PORT MAP(PP_IN(3)(40), PP_IN(4)(40), HA_lev6_col40_inst1_port_S, HA_lev6_col40_inst1_port_COUT);
FA_lev6_col41_inst0: FA PORT MAP(PP_IN(0)(41), PP_IN(1)(41), PP_IN(2)(41), FA_lev6_col41_inst0_port_S, FA_lev6_col41_inst0_port_COUT);
HA_lev6_col42_inst0: HA PORT MAP(PP_IN(0)(42), PP_IN(1)(42), HA_lev6_col42_inst0_port_S, HA_lev6_col42_inst0_port_COUT);

-- Level no 6
HA_lev5_col16_inst0: HA PORT MAP(PP_IN(0)(16), PP_IN(1)(16), HA_lev5_col16_inst0_port_S, HA_lev5_col16_inst0_port_COUT);
HA_lev5_col17_inst0: HA PORT MAP(PP_IN(0)(17), PP_IN(1)(17), HA_lev5_col17_inst0_port_S, HA_lev5_col17_inst0_port_COUT);
FA_lev5_col18_inst0: FA PORT MAP(PP_IN(0)(18), PP_IN(1)(18), PP_IN(2)(18), FA_lev5_col18_inst0_port_S, FA_lev5_col18_inst0_port_COUT);
HA_lev5_col18_inst1: HA PORT MAP(PP_IN(3)(18), PP_IN(4)(18), HA_lev5_col18_inst1_port_S, HA_lev5_col18_inst1_port_COUT);
FA_lev5_col19_inst0: FA PORT MAP(PP_IN(0)(19), PP_IN(1)(19), PP_IN(2)(19), FA_lev5_col19_inst0_port_S, FA_lev5_col19_inst0_port_COUT);
HA_lev5_col19_inst1: HA PORT MAP(PP_IN(3)(19), PP_IN(4)(19), HA_lev5_col19_inst1_port_S, HA_lev5_col19_inst1_port_COUT);
FA_lev5_col20_inst0: FA PORT MAP(PP_IN(0)(20), PP_IN(1)(20), PP_IN(2)(20), FA_lev5_col20_inst0_port_S, FA_lev5_col20_inst0_port_COUT);
FA_lev5_col20_inst1: FA PORT MAP(PP_IN(3)(20), PP_IN(4)(20), PP_IN(5)(20), FA_lev5_col20_inst1_port_S, FA_lev5_col20_inst1_port_COUT);
HA_lev5_col20_inst2: HA PORT MAP(PP_IN(6)(20), PP_IN(7)(20), HA_lev5_col20_inst2_port_S, HA_lev5_col20_inst2_port_COUT);
FA_lev5_col21_inst0: FA PORT MAP(PP_IN(0)(21), PP_IN(1)(21), PP_IN(2)(21), FA_lev5_col21_inst0_port_S, FA_lev5_col21_inst0_port_COUT);
FA_lev5_col21_inst1: FA PORT MAP(PP_IN(3)(21), PP_IN(4)(21), PP_IN(5)(21), FA_lev5_col21_inst1_port_S, FA_lev5_col21_inst1_port_COUT);
HA_lev5_col21_inst2: HA PORT MAP(PP_IN(6)(21), PP_IN(7)(21), HA_lev5_col21_inst2_port_S, HA_lev5_col21_inst2_port_COUT);
FA_lev5_col22_inst0: FA PORT MAP(PP_IN(0)(22), PP_IN(1)(22), PP_IN(2)(22), FA_lev5_col22_inst0_port_S, FA_lev5_col22_inst0_port_COUT);
FA_lev5_col22_inst1: FA PORT MAP(PP_IN(3)(22), PP_IN(4)(22), PP_IN(5)(22), FA_lev5_col22_inst1_port_S, FA_lev5_col22_inst1_port_COUT);
FA_lev5_col22_inst2: FA PORT MAP(PP_IN(6)(22), PP_IN(7)(22), PP_IN(8)(22), FA_lev5_col22_inst2_port_S, FA_lev5_col22_inst2_port_COUT);
HA_lev5_col22_inst3: HA PORT MAP(PP_IN(9)(22), PP_IN(10)(22), HA_lev5_col22_inst3_port_S, HA_lev5_col22_inst3_port_COUT);
FA_lev5_col23_inst0: FA PORT MAP(PP_IN(0)(23), PP_IN(1)(23), PP_IN(2)(23), FA_lev5_col23_inst0_port_S, FA_lev5_col23_inst0_port_COUT);
FA_lev5_col23_inst1: FA PORT MAP(PP_IN(3)(23), PP_IN(4)(23), PP_IN(5)(23), FA_lev5_col23_inst1_port_S, FA_lev5_col23_inst1_port_COUT);
FA_lev5_col23_inst2: FA PORT MAP(PP_IN(6)(23), PP_IN(7)(23), PP_IN(8)(23), FA_lev5_col23_inst2_port_S, FA_lev5_col23_inst2_port_COUT);
HA_lev5_col23_inst3: HA PORT MAP(PP_IN(9)(23), PP_IN(10)(23), HA_lev5_col23_inst3_port_S, HA_lev5_col23_inst3_port_COUT);
FA_lev5_col24_inst0: FA PORT MAP(HA_lev6_col24_inst0_port_S, PP_IN(2)(24), PP_IN(3)(24), FA_lev5_col24_inst0_port_S, FA_lev5_col24_inst0_port_COUT);
FA_lev5_col24_inst1: FA PORT MAP(PP_IN(4)(24), PP_IN(5)(24), PP_IN(6)(24), FA_lev5_col24_inst1_port_S, FA_lev5_col24_inst1_port_COUT);
FA_lev5_col24_inst2: FA PORT MAP(PP_IN(7)(24), PP_IN(8)(24), PP_IN(9)(24), FA_lev5_col24_inst2_port_S, FA_lev5_col24_inst2_port_COUT);
FA_lev5_col24_inst3: FA PORT MAP(PP_IN(10)(24), PP_IN(11)(24), PP_IN(12)(24), FA_lev5_col24_inst3_port_S, FA_lev5_col24_inst3_port_COUT);
FA_lev5_col25_inst0: FA PORT MAP(HA_lev6_col25_inst0_port_S, PP_IN(2)(25), PP_IN(3)(25), FA_lev5_col25_inst0_port_S, FA_lev5_col25_inst0_port_COUT);
FA_lev5_col25_inst1: FA PORT MAP(PP_IN(4)(25), PP_IN(5)(25), PP_IN(6)(25), FA_lev5_col25_inst1_port_S, FA_lev5_col25_inst1_port_COUT);
FA_lev5_col25_inst2: FA PORT MAP(PP_IN(7)(25), PP_IN(8)(25), PP_IN(9)(25), FA_lev5_col25_inst2_port_S, FA_lev5_col25_inst2_port_COUT);
FA_lev5_col25_inst3: FA PORT MAP(PP_IN(10)(25), PP_IN(11)(25), PP_IN(12)(25), FA_lev5_col25_inst3_port_S, FA_lev5_col25_inst3_port_COUT);
FA_lev5_col26_inst0: FA PORT MAP(FA_lev6_col26_inst0_port_S, HA_lev6_col26_inst1_port_S, PP_IN(5)(26), FA_lev5_col26_inst0_port_S, FA_lev5_col26_inst0_port_COUT);
FA_lev5_col26_inst1: FA PORT MAP(PP_IN(6)(26), PP_IN(7)(26), PP_IN(8)(26), FA_lev5_col26_inst1_port_S, FA_lev5_col26_inst1_port_COUT);
FA_lev5_col26_inst2: FA PORT MAP(PP_IN(9)(26), PP_IN(10)(26), PP_IN(11)(26), FA_lev5_col26_inst2_port_S, FA_lev5_col26_inst2_port_COUT);
FA_lev5_col26_inst3: FA PORT MAP(PP_IN(12)(26), PP_IN(13)(26), PP_IN(14)(26), FA_lev5_col26_inst3_port_S, FA_lev5_col26_inst3_port_COUT);
FA_lev5_col27_inst0: FA PORT MAP(FA_lev6_col27_inst0_port_S, HA_lev6_col27_inst1_port_S, PP_IN(5)(27), FA_lev5_col27_inst0_port_S, FA_lev5_col27_inst0_port_COUT);
FA_lev5_col27_inst1: FA PORT MAP(PP_IN(6)(27), PP_IN(7)(27), PP_IN(8)(27), FA_lev5_col27_inst1_port_S, FA_lev5_col27_inst1_port_COUT);
FA_lev5_col27_inst2: FA PORT MAP(PP_IN(9)(27), PP_IN(10)(27), PP_IN(11)(27), FA_lev5_col27_inst2_port_S, FA_lev5_col27_inst2_port_COUT);
FA_lev5_col27_inst3: FA PORT MAP(PP_IN(12)(27), PP_IN(13)(27), FA_lev6_col26_inst0_port_COUT, FA_lev5_col27_inst3_port_S, FA_lev5_col27_inst3_port_COUT);
FA_lev5_col28_inst0: FA PORT MAP(FA_lev6_col28_inst0_port_S, FA_lev6_col28_inst1_port_S, HA_lev6_col28_inst2_port_S, FA_lev5_col28_inst0_port_S, FA_lev5_col28_inst0_port_COUT);
FA_lev5_col28_inst1: FA PORT MAP(PP_IN(8)(28), PP_IN(9)(28), PP_IN(10)(28), FA_lev5_col28_inst1_port_S, FA_lev5_col28_inst1_port_COUT);
FA_lev5_col28_inst2: FA PORT MAP(PP_IN(11)(28), PP_IN(12)(28), PP_IN(13)(28), FA_lev5_col28_inst2_port_S, FA_lev5_col28_inst2_port_COUT);
FA_lev5_col28_inst3: FA PORT MAP(PP_IN(14)(28), PP_IN(15)(28), FA_lev6_col27_inst0_port_COUT, FA_lev5_col28_inst3_port_S, FA_lev5_col28_inst3_port_COUT);
FA_lev5_col29_inst0: FA PORT MAP(FA_lev6_col29_inst0_port_S, FA_lev6_col29_inst1_port_S, HA_lev6_col29_inst2_port_S, FA_lev5_col29_inst0_port_S, FA_lev5_col29_inst0_port_COUT);
FA_lev5_col29_inst1: FA PORT MAP(PP_IN(8)(29), PP_IN(9)(29), PP_IN(10)(29), FA_lev5_col29_inst1_port_S, FA_lev5_col29_inst1_port_COUT);
FA_lev5_col29_inst2: FA PORT MAP(PP_IN(11)(29), PP_IN(12)(29), PP_IN(13)(29), FA_lev5_col29_inst2_port_S, FA_lev5_col29_inst2_port_COUT);
FA_lev5_col29_inst3: FA PORT MAP(PP_IN(14)(29), FA_lev6_col28_inst0_port_COUT, FA_lev6_col28_inst1_port_COUT, FA_lev5_col29_inst3_port_S, FA_lev5_col29_inst3_port_COUT);
FA_lev5_col30_inst0: FA PORT MAP(FA_lev6_col30_inst0_port_S, FA_lev6_col30_inst1_port_S, FA_lev6_col30_inst2_port_S, FA_lev5_col30_inst0_port_S, FA_lev5_col30_inst0_port_COUT);
FA_lev5_col30_inst1: FA PORT MAP(HA_lev6_col30_inst3_port_S, PP_IN(11)(30), PP_IN(12)(30), FA_lev5_col30_inst1_port_S, FA_lev5_col30_inst1_port_COUT);
FA_lev5_col30_inst2: FA PORT MAP(PP_IN(13)(30), PP_IN(14)(30), PP_IN(15)(30), FA_lev5_col30_inst2_port_S, FA_lev5_col30_inst2_port_COUT);
FA_lev5_col30_inst3: FA PORT MAP(PP_IN(16)(30), FA_lev6_col29_inst0_port_COUT, FA_lev6_col29_inst1_port_COUT, FA_lev5_col30_inst3_port_S, FA_lev5_col30_inst3_port_COUT);
FA_lev5_col31_inst0: FA PORT MAP(FA_lev6_col31_inst0_port_S, FA_lev6_col31_inst1_port_S, FA_lev6_col31_inst2_port_S, FA_lev5_col31_inst0_port_S, FA_lev5_col31_inst0_port_COUT);
FA_lev5_col31_inst1: FA PORT MAP(HA_lev6_col31_inst3_port_S, PP_IN(11)(31), PP_IN(12)(31), FA_lev5_col31_inst1_port_S, FA_lev5_col31_inst1_port_COUT);
FA_lev5_col31_inst2: FA PORT MAP(PP_IN(13)(31), PP_IN(14)(31), PP_IN(15)(31), FA_lev5_col31_inst2_port_S, FA_lev5_col31_inst2_port_COUT);
FA_lev5_col31_inst3: FA PORT MAP(FA_lev6_col30_inst0_port_COUT, FA_lev6_col30_inst1_port_COUT, FA_lev6_col30_inst2_port_COUT, FA_lev5_col31_inst3_port_S, FA_lev5_col31_inst3_port_COUT);
FA_lev5_col32_inst0: FA PORT MAP(FA_lev6_col32_inst0_port_S, FA_lev6_col32_inst1_port_S, FA_lev6_col32_inst2_port_S, FA_lev5_col32_inst0_port_S, FA_lev5_col32_inst0_port_COUT);
FA_lev5_col32_inst1: FA PORT MAP(FA_lev6_col32_inst3_port_S, PP_IN(12)(32), PP_IN(13)(32), FA_lev5_col32_inst1_port_S, FA_lev5_col32_inst1_port_COUT);
FA_lev5_col32_inst2: FA PORT MAP(PP_IN(14)(32), PP_IN(15)(32), PP_IN(16)(32), FA_lev5_col32_inst2_port_S, FA_lev5_col32_inst2_port_COUT);
FA_lev5_col32_inst3: FA PORT MAP(FA_lev6_col31_inst0_port_COUT, FA_lev6_col31_inst1_port_COUT, FA_lev6_col31_inst2_port_COUT, FA_lev5_col32_inst3_port_S, FA_lev5_col32_inst3_port_COUT);
FA_lev5_col33_inst0: FA PORT MAP(FA_lev6_col33_inst0_port_S, FA_lev6_col33_inst1_port_S, FA_lev6_col33_inst2_port_S, FA_lev5_col33_inst0_port_S, FA_lev5_col33_inst0_port_COUT);
FA_lev5_col33_inst1: FA PORT MAP(FA_lev6_col33_inst3_port_S, PP_IN(12)(33), PP_IN(13)(33), FA_lev5_col33_inst1_port_S, FA_lev5_col33_inst1_port_COUT);
FA_lev5_col33_inst2: FA PORT MAP(PP_IN(14)(33), PP_IN(15)(33), PP_IN(16)(33), FA_lev5_col33_inst2_port_S, FA_lev5_col33_inst2_port_COUT);
FA_lev5_col33_inst3: FA PORT MAP(FA_lev6_col32_inst0_port_COUT, FA_lev6_col32_inst1_port_COUT, FA_lev6_col32_inst2_port_COUT, FA_lev5_col33_inst3_port_S, FA_lev5_col33_inst3_port_COUT);
FA_lev5_col34_inst0: FA PORT MAP(FA_lev6_col34_inst0_port_S, FA_lev6_col34_inst1_port_S, FA_lev6_col34_inst2_port_S, FA_lev5_col34_inst0_port_S, FA_lev5_col34_inst0_port_COUT);
FA_lev5_col34_inst1: FA PORT MAP(FA_lev6_col34_inst3_port_S, PP_IN(12)(34), PP_IN(13)(34), FA_lev5_col34_inst1_port_S, FA_lev5_col34_inst1_port_COUT);
FA_lev5_col34_inst2: FA PORT MAP(PP_IN(14)(34), PP_IN(15)(34), PP_IN(16)(34), FA_lev5_col34_inst2_port_S, FA_lev5_col34_inst2_port_COUT);
FA_lev5_col34_inst3: FA PORT MAP(FA_lev6_col33_inst0_port_COUT, FA_lev6_col33_inst1_port_COUT, FA_lev6_col33_inst2_port_COUT, FA_lev5_col34_inst3_port_S, FA_lev5_col34_inst3_port_COUT);
FA_lev5_col35_inst0: FA PORT MAP(FA_lev6_col35_inst0_port_S, FA_lev6_col35_inst1_port_S, FA_lev6_col35_inst2_port_S, FA_lev5_col35_inst0_port_S, FA_lev5_col35_inst0_port_COUT);
FA_lev5_col35_inst1: FA PORT MAP(FA_lev6_col35_inst3_port_S, PP_IN(12)(35), PP_IN(13)(35), FA_lev5_col35_inst1_port_S, FA_lev5_col35_inst1_port_COUT);
FA_lev5_col35_inst2: FA PORT MAP(PP_IN(14)(35), PP_IN(15)(35), PP_IN(16)(35), FA_lev5_col35_inst2_port_S, FA_lev5_col35_inst2_port_COUT);
FA_lev5_col35_inst3: FA PORT MAP(FA_lev6_col34_inst0_port_COUT, FA_lev6_col34_inst1_port_COUT, FA_lev6_col34_inst2_port_COUT, FA_lev5_col35_inst3_port_S, FA_lev5_col35_inst3_port_COUT);
FA_lev5_col36_inst0: FA PORT MAP(FA_lev6_col36_inst0_port_S, FA_lev6_col36_inst1_port_S, FA_lev6_col36_inst2_port_S, FA_lev5_col36_inst0_port_S, FA_lev5_col36_inst0_port_COUT);
FA_lev5_col36_inst1: FA PORT MAP(HA_lev6_col36_inst3_port_S, PP_IN(11)(36), PP_IN(12)(36), FA_lev5_col36_inst1_port_S, FA_lev5_col36_inst1_port_COUT);
FA_lev5_col36_inst2: FA PORT MAP(PP_IN(13)(36), PP_IN(14)(36), PP_IN(15)(36), FA_lev5_col36_inst2_port_S, FA_lev5_col36_inst2_port_COUT);
FA_lev5_col36_inst3: FA PORT MAP(FA_lev6_col35_inst0_port_COUT, FA_lev6_col35_inst1_port_COUT, FA_lev6_col35_inst2_port_COUT, FA_lev5_col36_inst3_port_S, FA_lev5_col36_inst3_port_COUT);
FA_lev5_col37_inst0: FA PORT MAP(FA_lev6_col37_inst0_port_S, FA_lev6_col37_inst1_port_S, FA_lev6_col37_inst2_port_S, FA_lev5_col37_inst0_port_S, FA_lev5_col37_inst0_port_COUT);
FA_lev5_col37_inst1: FA PORT MAP(PP_IN(9)(37), PP_IN(10)(37), PP_IN(11)(37), FA_lev5_col37_inst1_port_S, FA_lev5_col37_inst1_port_COUT);
FA_lev5_col37_inst2: FA PORT MAP(PP_IN(12)(37), PP_IN(13)(37), PP_IN(14)(37), FA_lev5_col37_inst2_port_S, FA_lev5_col37_inst2_port_COUT);
FA_lev5_col37_inst3: FA PORT MAP(FA_lev6_col36_inst0_port_COUT, FA_lev6_col36_inst1_port_COUT, FA_lev6_col36_inst2_port_COUT, FA_lev5_col37_inst3_port_S, FA_lev5_col37_inst3_port_COUT);
FA_lev5_col38_inst0: FA PORT MAP(FA_lev6_col38_inst0_port_S, FA_lev6_col38_inst1_port_S, HA_lev6_col38_inst2_port_S, FA_lev5_col38_inst0_port_S, FA_lev5_col38_inst0_port_COUT);
FA_lev5_col38_inst1: FA PORT MAP(PP_IN(8)(38), PP_IN(9)(38), PP_IN(10)(38), FA_lev5_col38_inst1_port_S, FA_lev5_col38_inst1_port_COUT);
FA_lev5_col38_inst2: FA PORT MAP(PP_IN(11)(38), PP_IN(12)(38), PP_IN(13)(38), FA_lev5_col38_inst2_port_S, FA_lev5_col38_inst2_port_COUT);
FA_lev5_col38_inst3: FA PORT MAP(PP_IN(14)(38), FA_lev6_col37_inst0_port_COUT, FA_lev6_col37_inst1_port_COUT, FA_lev5_col38_inst3_port_S, FA_lev5_col38_inst3_port_COUT);
FA_lev5_col39_inst0: FA PORT MAP(FA_lev6_col39_inst0_port_S, FA_lev6_col39_inst1_port_S, PP_IN(6)(39), FA_lev5_col39_inst0_port_S, FA_lev5_col39_inst0_port_COUT);
FA_lev5_col39_inst1: FA PORT MAP(PP_IN(7)(39), PP_IN(8)(39), PP_IN(9)(39), FA_lev5_col39_inst1_port_S, FA_lev5_col39_inst1_port_COUT);
FA_lev5_col39_inst2: FA PORT MAP(PP_IN(10)(39), PP_IN(11)(39), PP_IN(12)(39), FA_lev5_col39_inst2_port_S, FA_lev5_col39_inst2_port_COUT);
FA_lev5_col39_inst3: FA PORT MAP(PP_IN(13)(39), FA_lev6_col38_inst0_port_COUT, FA_lev6_col38_inst1_port_COUT, FA_lev5_col39_inst3_port_S, FA_lev5_col39_inst3_port_COUT);
FA_lev5_col40_inst0: FA PORT MAP(FA_lev6_col40_inst0_port_S, HA_lev6_col40_inst1_port_S, PP_IN(5)(40), FA_lev5_col40_inst0_port_S, FA_lev5_col40_inst0_port_COUT);
FA_lev5_col40_inst1: FA PORT MAP(PP_IN(6)(40), PP_IN(7)(40), PP_IN(8)(40), FA_lev5_col40_inst1_port_S, FA_lev5_col40_inst1_port_COUT);
FA_lev5_col40_inst2: FA PORT MAP(PP_IN(9)(40), PP_IN(10)(40), PP_IN(11)(40), FA_lev5_col40_inst2_port_S, FA_lev5_col40_inst2_port_COUT);
FA_lev5_col40_inst3: FA PORT MAP(PP_IN(12)(40), PP_IN(13)(40), FA_lev6_col39_inst0_port_COUT, FA_lev5_col40_inst3_port_S, FA_lev5_col40_inst3_port_COUT);
FA_lev5_col41_inst0: FA PORT MAP(FA_lev6_col41_inst0_port_S, PP_IN(3)(41), PP_IN(4)(41), FA_lev5_col41_inst0_port_S, FA_lev5_col41_inst0_port_COUT);
FA_lev5_col41_inst1: FA PORT MAP(PP_IN(5)(41), PP_IN(6)(41), PP_IN(7)(41), FA_lev5_col41_inst1_port_S, FA_lev5_col41_inst1_port_COUT);
FA_lev5_col41_inst2: FA PORT MAP(PP_IN(8)(41), PP_IN(9)(41), PP_IN(10)(41), FA_lev5_col41_inst2_port_S, FA_lev5_col41_inst2_port_COUT);
FA_lev5_col41_inst3: FA PORT MAP(PP_IN(11)(41), PP_IN(12)(41), FA_lev6_col40_inst0_port_COUT, FA_lev5_col41_inst3_port_S, FA_lev5_col41_inst3_port_COUT);
FA_lev5_col42_inst0: FA PORT MAP(HA_lev6_col42_inst0_port_S, PP_IN(2)(42), PP_IN(3)(42), FA_lev5_col42_inst0_port_S, FA_lev5_col42_inst0_port_COUT);
FA_lev5_col42_inst1: FA PORT MAP(PP_IN(4)(42), PP_IN(5)(42), PP_IN(6)(42), FA_lev5_col42_inst1_port_S, FA_lev5_col42_inst1_port_COUT);
FA_lev5_col42_inst2: FA PORT MAP(PP_IN(7)(42), PP_IN(8)(42), PP_IN(9)(42), FA_lev5_col42_inst2_port_S, FA_lev5_col42_inst2_port_COUT);
FA_lev5_col42_inst3: FA PORT MAP(PP_IN(10)(42), PP_IN(11)(42), PP_IN(12)(42), FA_lev5_col42_inst3_port_S, FA_lev5_col42_inst3_port_COUT);
FA_lev5_col43_inst0: FA PORT MAP(PP_IN(0)(43), PP_IN(1)(43), PP_IN(2)(43), FA_lev5_col43_inst0_port_S, FA_lev5_col43_inst0_port_COUT);
FA_lev5_col43_inst1: FA PORT MAP(PP_IN(3)(43), PP_IN(4)(43), PP_IN(5)(43), FA_lev5_col43_inst1_port_S, FA_lev5_col43_inst1_port_COUT);
FA_lev5_col43_inst2: FA PORT MAP(PP_IN(6)(43), PP_IN(7)(43), PP_IN(8)(43), FA_lev5_col43_inst2_port_S, FA_lev5_col43_inst2_port_COUT);
FA_lev5_col43_inst3: FA PORT MAP(PP_IN(9)(43), PP_IN(10)(43), PP_IN(11)(43), FA_lev5_col43_inst3_port_S, FA_lev5_col43_inst3_port_COUT);
FA_lev5_col44_inst0: FA PORT MAP(PP_IN(0)(44), PP_IN(1)(44), PP_IN(2)(44), FA_lev5_col44_inst0_port_S, FA_lev5_col44_inst0_port_COUT);
FA_lev5_col44_inst1: FA PORT MAP(PP_IN(3)(44), PP_IN(4)(44), PP_IN(5)(44), FA_lev5_col44_inst1_port_S, FA_lev5_col44_inst1_port_COUT);
FA_lev5_col44_inst2: FA PORT MAP(PP_IN(6)(44), PP_IN(7)(44), PP_IN(8)(44), FA_lev5_col44_inst2_port_S, FA_lev5_col44_inst2_port_COUT);
HA_lev5_col44_inst3: HA PORT MAP(PP_IN(9)(44), PP_IN(10)(44), HA_lev5_col44_inst3_port_S, HA_lev5_col44_inst3_port_COUT);
FA_lev5_col45_inst0: FA PORT MAP(PP_IN(0)(45), PP_IN(1)(45), PP_IN(2)(45), FA_lev5_col45_inst0_port_S, FA_lev5_col45_inst0_port_COUT);
FA_lev5_col45_inst1: FA PORT MAP(PP_IN(3)(45), PP_IN(4)(45), PP_IN(5)(45), FA_lev5_col45_inst1_port_S, FA_lev5_col45_inst1_port_COUT);
FA_lev5_col45_inst2: FA PORT MAP(PP_IN(6)(45), PP_IN(7)(45), PP_IN(8)(45), FA_lev5_col45_inst2_port_S, FA_lev5_col45_inst2_port_COUT);
FA_lev5_col46_inst0: FA PORT MAP(PP_IN(0)(46), PP_IN(1)(46), PP_IN(2)(46), FA_lev5_col46_inst0_port_S, FA_lev5_col46_inst0_port_COUT);
FA_lev5_col46_inst1: FA PORT MAP(PP_IN(3)(46), PP_IN(4)(46), PP_IN(5)(46), FA_lev5_col46_inst1_port_S, FA_lev5_col46_inst1_port_COUT);
HA_lev5_col46_inst2: HA PORT MAP(PP_IN(6)(46), PP_IN(7)(46), HA_lev5_col46_inst2_port_S, HA_lev5_col46_inst2_port_COUT);
FA_lev5_col47_inst0: FA PORT MAP(PP_IN(0)(47), PP_IN(1)(47), PP_IN(2)(47), FA_lev5_col47_inst0_port_S, FA_lev5_col47_inst0_port_COUT);
FA_lev5_col47_inst1: FA PORT MAP(PP_IN(3)(47), PP_IN(4)(47), PP_IN(5)(47), FA_lev5_col47_inst1_port_S, FA_lev5_col47_inst1_port_COUT);
FA_lev5_col48_inst0: FA PORT MAP(PP_IN(0)(48), PP_IN(1)(48), PP_IN(2)(48), FA_lev5_col48_inst0_port_S, FA_lev5_col48_inst0_port_COUT);
HA_lev5_col48_inst1: HA PORT MAP(PP_IN(3)(48), PP_IN(4)(48), HA_lev5_col48_inst1_port_S, HA_lev5_col48_inst1_port_COUT);
FA_lev5_col49_inst0: FA PORT MAP(PP_IN(0)(49), PP_IN(1)(49), PP_IN(2)(49), FA_lev5_col49_inst0_port_S, FA_lev5_col49_inst0_port_COUT);
HA_lev5_col50_inst0: HA PORT MAP(PP_IN(0)(50), PP_IN(1)(50), HA_lev5_col50_inst0_port_S, HA_lev5_col50_inst0_port_COUT);

-- Level no 5
HA_lev4_col10_inst0: HA PORT MAP(PP_IN(0)(10), PP_IN(1)(10), HA_lev4_col10_inst0_port_S, HA_lev4_col10_inst0_port_COUT);
HA_lev4_col11_inst0: HA PORT MAP(PP_IN(0)(11), PP_IN(1)(11), HA_lev4_col11_inst0_port_S, HA_lev4_col11_inst0_port_COUT);
FA_lev4_col12_inst0: FA PORT MAP(PP_IN(0)(12), PP_IN(1)(12), PP_IN(2)(12), FA_lev4_col12_inst0_port_S, FA_lev4_col12_inst0_port_COUT);
HA_lev4_col12_inst1: HA PORT MAP(PP_IN(3)(12), PP_IN(4)(12), HA_lev4_col12_inst1_port_S, HA_lev4_col12_inst1_port_COUT);
FA_lev4_col13_inst0: FA PORT MAP(PP_IN(0)(13), PP_IN(1)(13), PP_IN(2)(13), FA_lev4_col13_inst0_port_S, FA_lev4_col13_inst0_port_COUT);
HA_lev4_col13_inst1: HA PORT MAP(PP_IN(3)(13), PP_IN(4)(13), HA_lev4_col13_inst1_port_S, HA_lev4_col13_inst1_port_COUT);
FA_lev4_col14_inst0: FA PORT MAP(PP_IN(0)(14), PP_IN(1)(14), PP_IN(2)(14), FA_lev4_col14_inst0_port_S, FA_lev4_col14_inst0_port_COUT);
FA_lev4_col14_inst1: FA PORT MAP(PP_IN(3)(14), PP_IN(4)(14), PP_IN(5)(14), FA_lev4_col14_inst1_port_S, FA_lev4_col14_inst1_port_COUT);
HA_lev4_col14_inst2: HA PORT MAP(PP_IN(6)(14), PP_IN(7)(14), HA_lev4_col14_inst2_port_S, HA_lev4_col14_inst2_port_COUT);
FA_lev4_col15_inst0: FA PORT MAP(PP_IN(0)(15), PP_IN(1)(15), PP_IN(2)(15), FA_lev4_col15_inst0_port_S, FA_lev4_col15_inst0_port_COUT);
FA_lev4_col15_inst1: FA PORT MAP(PP_IN(3)(15), PP_IN(4)(15), PP_IN(5)(15), FA_lev4_col15_inst1_port_S, FA_lev4_col15_inst1_port_COUT);
HA_lev4_col15_inst2: HA PORT MAP(PP_IN(6)(15), PP_IN(7)(15), HA_lev4_col15_inst2_port_S, HA_lev4_col15_inst2_port_COUT);
FA_lev4_col16_inst0: FA PORT MAP(HA_lev5_col16_inst0_port_S, PP_IN(2)(16), PP_IN(3)(16), FA_lev4_col16_inst0_port_S, FA_lev4_col16_inst0_port_COUT);
FA_lev4_col16_inst1: FA PORT MAP(PP_IN(4)(16), PP_IN(5)(16), PP_IN(6)(16), FA_lev4_col16_inst1_port_S, FA_lev4_col16_inst1_port_COUT);
FA_lev4_col16_inst2: FA PORT MAP(PP_IN(7)(16), PP_IN(8)(16), PP_IN(9)(16), FA_lev4_col16_inst2_port_S, FA_lev4_col16_inst2_port_COUT);
FA_lev4_col17_inst0: FA PORT MAP(HA_lev5_col17_inst0_port_S, PP_IN(2)(17), PP_IN(3)(17), FA_lev4_col17_inst0_port_S, FA_lev4_col17_inst0_port_COUT);
FA_lev4_col17_inst1: FA PORT MAP(PP_IN(4)(17), PP_IN(5)(17), PP_IN(6)(17), FA_lev4_col17_inst1_port_S, FA_lev4_col17_inst1_port_COUT);
FA_lev4_col17_inst2: FA PORT MAP(PP_IN(7)(17), PP_IN(8)(17), HA_lev5_col16_inst0_port_COUT, FA_lev4_col17_inst2_port_S, FA_lev4_col17_inst2_port_COUT);
FA_lev4_col18_inst0: FA PORT MAP(FA_lev5_col18_inst0_port_S, HA_lev5_col18_inst1_port_S, PP_IN(5)(18), FA_lev4_col18_inst0_port_S, FA_lev4_col18_inst0_port_COUT);
FA_lev4_col18_inst1: FA PORT MAP(PP_IN(6)(18), PP_IN(7)(18), PP_IN(8)(18), FA_lev4_col18_inst1_port_S, FA_lev4_col18_inst1_port_COUT);
FA_lev4_col18_inst2: FA PORT MAP(PP_IN(9)(18), PP_IN(10)(18), HA_lev5_col17_inst0_port_COUT, FA_lev4_col18_inst2_port_S, FA_lev4_col18_inst2_port_COUT);
FA_lev4_col19_inst0: FA PORT MAP(FA_lev5_col19_inst0_port_S, HA_lev5_col19_inst1_port_S, PP_IN(5)(19), FA_lev4_col19_inst0_port_S, FA_lev4_col19_inst0_port_COUT);
FA_lev4_col19_inst1: FA PORT MAP(PP_IN(6)(19), PP_IN(7)(19), PP_IN(8)(19), FA_lev4_col19_inst1_port_S, FA_lev4_col19_inst1_port_COUT);
FA_lev4_col19_inst2: FA PORT MAP(PP_IN(9)(19), FA_lev5_col18_inst0_port_COUT, HA_lev5_col18_inst1_port_COUT, FA_lev4_col19_inst2_port_S, FA_lev4_col19_inst2_port_COUT);
FA_lev4_col20_inst0: FA PORT MAP(FA_lev5_col20_inst0_port_S, FA_lev5_col20_inst1_port_S, HA_lev5_col20_inst2_port_S, FA_lev4_col20_inst0_port_S, FA_lev4_col20_inst0_port_COUT);
FA_lev4_col20_inst1: FA PORT MAP(PP_IN(8)(20), PP_IN(9)(20), PP_IN(10)(20), FA_lev4_col20_inst1_port_S, FA_lev4_col20_inst1_port_COUT);
FA_lev4_col20_inst2: FA PORT MAP(PP_IN(11)(20), FA_lev5_col19_inst0_port_COUT, HA_lev5_col19_inst1_port_COUT, FA_lev4_col20_inst2_port_S, FA_lev4_col20_inst2_port_COUT);
FA_lev4_col21_inst0: FA PORT MAP(FA_lev5_col21_inst0_port_S, FA_lev5_col21_inst1_port_S, HA_lev5_col21_inst2_port_S, FA_lev4_col21_inst0_port_S, FA_lev4_col21_inst0_port_COUT);
FA_lev4_col21_inst1: FA PORT MAP(PP_IN(8)(21), PP_IN(9)(21), PP_IN(10)(21), FA_lev4_col21_inst1_port_S, FA_lev4_col21_inst1_port_COUT);
FA_lev4_col21_inst2: FA PORT MAP(FA_lev5_col20_inst0_port_COUT, FA_lev5_col20_inst1_port_COUT, HA_lev5_col20_inst2_port_COUT, FA_lev4_col21_inst2_port_S, FA_lev4_col21_inst2_port_COUT);
FA_lev4_col22_inst0: FA PORT MAP(FA_lev5_col22_inst0_port_S, FA_lev5_col22_inst1_port_S, FA_lev5_col22_inst2_port_S, FA_lev4_col22_inst0_port_S, FA_lev4_col22_inst0_port_COUT);
FA_lev4_col22_inst1: FA PORT MAP(HA_lev5_col22_inst3_port_S, PP_IN(11)(22), PP_IN(12)(22), FA_lev4_col22_inst1_port_S, FA_lev4_col22_inst1_port_COUT);
FA_lev4_col22_inst2: FA PORT MAP(FA_lev5_col21_inst0_port_COUT, FA_lev5_col21_inst1_port_COUT, HA_lev5_col21_inst2_port_COUT, FA_lev4_col22_inst2_port_S, FA_lev4_col22_inst2_port_COUT);
FA_lev4_col23_inst0: FA PORT MAP(FA_lev5_col23_inst0_port_S, FA_lev5_col23_inst1_port_S, FA_lev5_col23_inst2_port_S, FA_lev4_col23_inst0_port_S, FA_lev4_col23_inst0_port_COUT);
FA_lev4_col23_inst1: FA PORT MAP(HA_lev5_col23_inst3_port_S, PP_IN(11)(23), FA_lev5_col22_inst0_port_COUT, FA_lev4_col23_inst1_port_S, FA_lev4_col23_inst1_port_COUT);
FA_lev4_col23_inst2: FA PORT MAP(FA_lev5_col22_inst1_port_COUT, FA_lev5_col22_inst2_port_COUT, HA_lev5_col22_inst3_port_COUT, FA_lev4_col23_inst2_port_S, FA_lev4_col23_inst2_port_COUT);
FA_lev4_col24_inst0: FA PORT MAP(FA_lev5_col24_inst0_port_S, FA_lev5_col24_inst1_port_S, FA_lev5_col24_inst2_port_S, FA_lev4_col24_inst0_port_S, FA_lev4_col24_inst0_port_COUT);
FA_lev4_col24_inst1: FA PORT MAP(FA_lev5_col24_inst3_port_S, PP_IN(13)(24), FA_lev5_col23_inst0_port_COUT, FA_lev4_col24_inst1_port_S, FA_lev4_col24_inst1_port_COUT);
FA_lev4_col24_inst2: FA PORT MAP(FA_lev5_col23_inst1_port_COUT, FA_lev5_col23_inst2_port_COUT, HA_lev5_col23_inst3_port_COUT, FA_lev4_col24_inst2_port_S, FA_lev4_col24_inst2_port_COUT);
FA_lev4_col25_inst0: FA PORT MAP(FA_lev5_col25_inst0_port_S, FA_lev5_col25_inst1_port_S, FA_lev5_col25_inst2_port_S, FA_lev4_col25_inst0_port_S, FA_lev4_col25_inst0_port_COUT);
FA_lev4_col25_inst1: FA PORT MAP(FA_lev5_col25_inst3_port_S, HA_lev6_col24_inst0_port_COUT, FA_lev5_col24_inst0_port_COUT, FA_lev4_col25_inst1_port_S, FA_lev4_col25_inst1_port_COUT);
FA_lev4_col25_inst2: FA PORT MAP(FA_lev5_col24_inst1_port_COUT, FA_lev5_col24_inst2_port_COUT, FA_lev5_col24_inst3_port_COUT, FA_lev4_col25_inst2_port_S, FA_lev4_col25_inst2_port_COUT);
FA_lev4_col26_inst0: FA PORT MAP(FA_lev5_col26_inst0_port_S, FA_lev5_col26_inst1_port_S, FA_lev5_col26_inst2_port_S, FA_lev4_col26_inst0_port_S, FA_lev4_col26_inst0_port_COUT);
FA_lev4_col26_inst1: FA PORT MAP(FA_lev5_col26_inst3_port_S, HA_lev6_col25_inst0_port_COUT, FA_lev5_col25_inst0_port_COUT, FA_lev4_col26_inst1_port_S, FA_lev4_col26_inst1_port_COUT);
FA_lev4_col26_inst2: FA PORT MAP(FA_lev5_col25_inst1_port_COUT, FA_lev5_col25_inst2_port_COUT, FA_lev5_col25_inst3_port_COUT, FA_lev4_col26_inst2_port_S, FA_lev4_col26_inst2_port_COUT);
FA_lev4_col27_inst0: FA PORT MAP(FA_lev5_col27_inst0_port_S, FA_lev5_col27_inst1_port_S, FA_lev5_col27_inst2_port_S, FA_lev4_col27_inst0_port_S, FA_lev4_col27_inst0_port_COUT);
FA_lev4_col27_inst1: FA PORT MAP(FA_lev5_col27_inst3_port_S, HA_lev6_col26_inst1_port_COUT, FA_lev5_col26_inst0_port_COUT, FA_lev4_col27_inst1_port_S, FA_lev4_col27_inst1_port_COUT);
FA_lev4_col27_inst2: FA PORT MAP(FA_lev5_col26_inst1_port_COUT, FA_lev5_col26_inst2_port_COUT, FA_lev5_col26_inst3_port_COUT, FA_lev4_col27_inst2_port_S, FA_lev4_col27_inst2_port_COUT);
FA_lev4_col28_inst0: FA PORT MAP(FA_lev5_col28_inst0_port_S, FA_lev5_col28_inst1_port_S, FA_lev5_col28_inst2_port_S, FA_lev4_col28_inst0_port_S, FA_lev4_col28_inst0_port_COUT);
FA_lev4_col28_inst1: FA PORT MAP(FA_lev5_col28_inst3_port_S, HA_lev6_col27_inst1_port_COUT, FA_lev5_col27_inst0_port_COUT, FA_lev4_col28_inst1_port_S, FA_lev4_col28_inst1_port_COUT);
FA_lev4_col28_inst2: FA PORT MAP(FA_lev5_col27_inst1_port_COUT, FA_lev5_col27_inst2_port_COUT, FA_lev5_col27_inst3_port_COUT, FA_lev4_col28_inst2_port_S, FA_lev4_col28_inst2_port_COUT);
FA_lev4_col29_inst0: FA PORT MAP(FA_lev5_col29_inst0_port_S, FA_lev5_col29_inst1_port_S, FA_lev5_col29_inst2_port_S, FA_lev4_col29_inst0_port_S, FA_lev4_col29_inst0_port_COUT);
FA_lev4_col29_inst1: FA PORT MAP(FA_lev5_col29_inst3_port_S, HA_lev6_col28_inst2_port_COUT, FA_lev5_col28_inst0_port_COUT, FA_lev4_col29_inst1_port_S, FA_lev4_col29_inst1_port_COUT);
FA_lev4_col29_inst2: FA PORT MAP(FA_lev5_col28_inst1_port_COUT, FA_lev5_col28_inst2_port_COUT, FA_lev5_col28_inst3_port_COUT, FA_lev4_col29_inst2_port_S, FA_lev4_col29_inst2_port_COUT);
FA_lev4_col30_inst0: FA PORT MAP(FA_lev5_col30_inst0_port_S, FA_lev5_col30_inst1_port_S, FA_lev5_col30_inst2_port_S, FA_lev4_col30_inst0_port_S, FA_lev4_col30_inst0_port_COUT);
FA_lev4_col30_inst1: FA PORT MAP(FA_lev5_col30_inst3_port_S, HA_lev6_col29_inst2_port_COUT, FA_lev5_col29_inst0_port_COUT, FA_lev4_col30_inst1_port_S, FA_lev4_col30_inst1_port_COUT);
FA_lev4_col30_inst2: FA PORT MAP(FA_lev5_col29_inst1_port_COUT, FA_lev5_col29_inst2_port_COUT, FA_lev5_col29_inst3_port_COUT, FA_lev4_col30_inst2_port_S, FA_lev4_col30_inst2_port_COUT);
FA_lev4_col31_inst0: FA PORT MAP(FA_lev5_col31_inst0_port_S, FA_lev5_col31_inst1_port_S, FA_lev5_col31_inst2_port_S, FA_lev4_col31_inst0_port_S, FA_lev4_col31_inst0_port_COUT);
FA_lev4_col31_inst1: FA PORT MAP(FA_lev5_col31_inst3_port_S, HA_lev6_col30_inst3_port_COUT, FA_lev5_col30_inst0_port_COUT, FA_lev4_col31_inst1_port_S, FA_lev4_col31_inst1_port_COUT);
FA_lev4_col31_inst2: FA PORT MAP(FA_lev5_col30_inst1_port_COUT, FA_lev5_col30_inst2_port_COUT, FA_lev5_col30_inst3_port_COUT, FA_lev4_col31_inst2_port_S, FA_lev4_col31_inst2_port_COUT);
FA_lev4_col32_inst0: FA PORT MAP(FA_lev5_col32_inst0_port_S, FA_lev5_col32_inst1_port_S, FA_lev5_col32_inst2_port_S, FA_lev4_col32_inst0_port_S, FA_lev4_col32_inst0_port_COUT);
FA_lev4_col32_inst1: FA PORT MAP(FA_lev5_col32_inst3_port_S, HA_lev6_col31_inst3_port_COUT, FA_lev5_col31_inst0_port_COUT, FA_lev4_col32_inst1_port_S, FA_lev4_col32_inst1_port_COUT);
FA_lev4_col32_inst2: FA PORT MAP(FA_lev5_col31_inst1_port_COUT, FA_lev5_col31_inst2_port_COUT, FA_lev5_col31_inst3_port_COUT, FA_lev4_col32_inst2_port_S, FA_lev4_col32_inst2_port_COUT);
FA_lev4_col33_inst0: FA PORT MAP(FA_lev5_col33_inst0_port_S, FA_lev5_col33_inst1_port_S, FA_lev5_col33_inst2_port_S, FA_lev4_col33_inst0_port_S, FA_lev4_col33_inst0_port_COUT);
FA_lev4_col33_inst1: FA PORT MAP(FA_lev5_col33_inst3_port_S, FA_lev6_col32_inst3_port_COUT, FA_lev5_col32_inst0_port_COUT, FA_lev4_col33_inst1_port_S, FA_lev4_col33_inst1_port_COUT);
FA_lev4_col33_inst2: FA PORT MAP(FA_lev5_col32_inst1_port_COUT, FA_lev5_col32_inst2_port_COUT, FA_lev5_col32_inst3_port_COUT, FA_lev4_col33_inst2_port_S, FA_lev4_col33_inst2_port_COUT);
FA_lev4_col34_inst0: FA PORT MAP(FA_lev5_col34_inst0_port_S, FA_lev5_col34_inst1_port_S, FA_lev5_col34_inst2_port_S, FA_lev4_col34_inst0_port_S, FA_lev4_col34_inst0_port_COUT);
FA_lev4_col34_inst1: FA PORT MAP(FA_lev5_col34_inst3_port_S, FA_lev6_col33_inst3_port_COUT, FA_lev5_col33_inst0_port_COUT, FA_lev4_col34_inst1_port_S, FA_lev4_col34_inst1_port_COUT);
FA_lev4_col34_inst2: FA PORT MAP(FA_lev5_col33_inst1_port_COUT, FA_lev5_col33_inst2_port_COUT, FA_lev5_col33_inst3_port_COUT, FA_lev4_col34_inst2_port_S, FA_lev4_col34_inst2_port_COUT);
FA_lev4_col35_inst0: FA PORT MAP(FA_lev5_col35_inst0_port_S, FA_lev5_col35_inst1_port_S, FA_lev5_col35_inst2_port_S, FA_lev4_col35_inst0_port_S, FA_lev4_col35_inst0_port_COUT);
FA_lev4_col35_inst1: FA PORT MAP(FA_lev5_col35_inst3_port_S, FA_lev6_col34_inst3_port_COUT, FA_lev5_col34_inst0_port_COUT, FA_lev4_col35_inst1_port_S, FA_lev4_col35_inst1_port_COUT);
FA_lev4_col35_inst2: FA PORT MAP(FA_lev5_col34_inst1_port_COUT, FA_lev5_col34_inst2_port_COUT, FA_lev5_col34_inst3_port_COUT, FA_lev4_col35_inst2_port_S, FA_lev4_col35_inst2_port_COUT);
FA_lev4_col36_inst0: FA PORT MAP(FA_lev5_col36_inst0_port_S, FA_lev5_col36_inst1_port_S, FA_lev5_col36_inst2_port_S, FA_lev4_col36_inst0_port_S, FA_lev4_col36_inst0_port_COUT);
FA_lev4_col36_inst1: FA PORT MAP(FA_lev5_col36_inst3_port_S, FA_lev6_col35_inst3_port_COUT, FA_lev5_col35_inst0_port_COUT, FA_lev4_col36_inst1_port_S, FA_lev4_col36_inst1_port_COUT);
FA_lev4_col36_inst2: FA PORT MAP(FA_lev5_col35_inst1_port_COUT, FA_lev5_col35_inst2_port_COUT, FA_lev5_col35_inst3_port_COUT, FA_lev4_col36_inst2_port_S, FA_lev4_col36_inst2_port_COUT);
FA_lev4_col37_inst0: FA PORT MAP(FA_lev5_col37_inst0_port_S, FA_lev5_col37_inst1_port_S, FA_lev5_col37_inst2_port_S, FA_lev4_col37_inst0_port_S, FA_lev4_col37_inst0_port_COUT);
FA_lev4_col37_inst1: FA PORT MAP(FA_lev5_col37_inst3_port_S, HA_lev6_col36_inst3_port_COUT, FA_lev5_col36_inst0_port_COUT, FA_lev4_col37_inst1_port_S, FA_lev4_col37_inst1_port_COUT);
FA_lev4_col37_inst2: FA PORT MAP(FA_lev5_col36_inst1_port_COUT, FA_lev5_col36_inst2_port_COUT, FA_lev5_col36_inst3_port_COUT, FA_lev4_col37_inst2_port_S, FA_lev4_col37_inst2_port_COUT);
FA_lev4_col38_inst0: FA PORT MAP(FA_lev5_col38_inst0_port_S, FA_lev5_col38_inst1_port_S, FA_lev5_col38_inst2_port_S, FA_lev4_col38_inst0_port_S, FA_lev4_col38_inst0_port_COUT);
FA_lev4_col38_inst1: FA PORT MAP(FA_lev5_col38_inst3_port_S, FA_lev6_col37_inst2_port_COUT, FA_lev5_col37_inst0_port_COUT, FA_lev4_col38_inst1_port_S, FA_lev4_col38_inst1_port_COUT);
FA_lev4_col38_inst2: FA PORT MAP(FA_lev5_col37_inst1_port_COUT, FA_lev5_col37_inst2_port_COUT, FA_lev5_col37_inst3_port_COUT, FA_lev4_col38_inst2_port_S, FA_lev4_col38_inst2_port_COUT);
FA_lev4_col39_inst0: FA PORT MAP(FA_lev5_col39_inst0_port_S, FA_lev5_col39_inst1_port_S, FA_lev5_col39_inst2_port_S, FA_lev4_col39_inst0_port_S, FA_lev4_col39_inst0_port_COUT);
FA_lev4_col39_inst1: FA PORT MAP(FA_lev5_col39_inst3_port_S, HA_lev6_col38_inst2_port_COUT, FA_lev5_col38_inst0_port_COUT, FA_lev4_col39_inst1_port_S, FA_lev4_col39_inst1_port_COUT);
FA_lev4_col39_inst2: FA PORT MAP(FA_lev5_col38_inst1_port_COUT, FA_lev5_col38_inst2_port_COUT, FA_lev5_col38_inst3_port_COUT, FA_lev4_col39_inst2_port_S, FA_lev4_col39_inst2_port_COUT);
FA_lev4_col40_inst0: FA PORT MAP(FA_lev5_col40_inst0_port_S, FA_lev5_col40_inst1_port_S, FA_lev5_col40_inst2_port_S, FA_lev4_col40_inst0_port_S, FA_lev4_col40_inst0_port_COUT);
FA_lev4_col40_inst1: FA PORT MAP(FA_lev5_col40_inst3_port_S, FA_lev6_col39_inst1_port_COUT, FA_lev5_col39_inst0_port_COUT, FA_lev4_col40_inst1_port_S, FA_lev4_col40_inst1_port_COUT);
FA_lev4_col40_inst2: FA PORT MAP(FA_lev5_col39_inst1_port_COUT, FA_lev5_col39_inst2_port_COUT, FA_lev5_col39_inst3_port_COUT, FA_lev4_col40_inst2_port_S, FA_lev4_col40_inst2_port_COUT);
FA_lev4_col41_inst0: FA PORT MAP(FA_lev5_col41_inst0_port_S, FA_lev5_col41_inst1_port_S, FA_lev5_col41_inst2_port_S, FA_lev4_col41_inst0_port_S, FA_lev4_col41_inst0_port_COUT);
FA_lev4_col41_inst1: FA PORT MAP(FA_lev5_col41_inst3_port_S, HA_lev6_col40_inst1_port_COUT, FA_lev5_col40_inst0_port_COUT, FA_lev4_col41_inst1_port_S, FA_lev4_col41_inst1_port_COUT);
FA_lev4_col41_inst2: FA PORT MAP(FA_lev5_col40_inst1_port_COUT, FA_lev5_col40_inst2_port_COUT, FA_lev5_col40_inst3_port_COUT, FA_lev4_col41_inst2_port_S, FA_lev4_col41_inst2_port_COUT);
FA_lev4_col42_inst0: FA PORT MAP(FA_lev5_col42_inst0_port_S, FA_lev5_col42_inst1_port_S, FA_lev5_col42_inst2_port_S, FA_lev4_col42_inst0_port_S, FA_lev4_col42_inst0_port_COUT);
FA_lev4_col42_inst1: FA PORT MAP(FA_lev5_col42_inst3_port_S, FA_lev6_col41_inst0_port_COUT, FA_lev5_col41_inst0_port_COUT, FA_lev4_col42_inst1_port_S, FA_lev4_col42_inst1_port_COUT);
FA_lev4_col42_inst2: FA PORT MAP(FA_lev5_col41_inst1_port_COUT, FA_lev5_col41_inst2_port_COUT, FA_lev5_col41_inst3_port_COUT, FA_lev4_col42_inst2_port_S, FA_lev4_col42_inst2_port_COUT);
FA_lev4_col43_inst0: FA PORT MAP(FA_lev5_col43_inst0_port_S, FA_lev5_col43_inst1_port_S, FA_lev5_col43_inst2_port_S, FA_lev4_col43_inst0_port_S, FA_lev4_col43_inst0_port_COUT);
FA_lev4_col43_inst1: FA PORT MAP(FA_lev5_col43_inst3_port_S, HA_lev6_col42_inst0_port_COUT, FA_lev5_col42_inst0_port_COUT, FA_lev4_col43_inst1_port_S, FA_lev4_col43_inst1_port_COUT);
FA_lev4_col43_inst2: FA PORT MAP(FA_lev5_col42_inst1_port_COUT, FA_lev5_col42_inst2_port_COUT, FA_lev5_col42_inst3_port_COUT, FA_lev4_col43_inst2_port_S, FA_lev4_col43_inst2_port_COUT);
FA_lev4_col44_inst0: FA PORT MAP(FA_lev5_col44_inst0_port_S, FA_lev5_col44_inst1_port_S, FA_lev5_col44_inst2_port_S, FA_lev4_col44_inst0_port_S, FA_lev4_col44_inst0_port_COUT);
FA_lev4_col44_inst1: FA PORT MAP(HA_lev5_col44_inst3_port_S, PP_IN(11)(44), FA_lev5_col43_inst0_port_COUT, FA_lev4_col44_inst1_port_S, FA_lev4_col44_inst1_port_COUT);
FA_lev4_col44_inst2: FA PORT MAP(FA_lev5_col43_inst1_port_COUT, FA_lev5_col43_inst2_port_COUT, FA_lev5_col43_inst3_port_COUT, FA_lev4_col44_inst2_port_S, FA_lev4_col44_inst2_port_COUT);
FA_lev4_col45_inst0: FA PORT MAP(FA_lev5_col45_inst0_port_S, FA_lev5_col45_inst1_port_S, FA_lev5_col45_inst2_port_S, FA_lev4_col45_inst0_port_S, FA_lev4_col45_inst0_port_COUT);
FA_lev4_col45_inst1: FA PORT MAP(PP_IN(9)(45), PP_IN(10)(45), FA_lev5_col44_inst0_port_COUT, FA_lev4_col45_inst1_port_S, FA_lev4_col45_inst1_port_COUT);
FA_lev4_col45_inst2: FA PORT MAP(FA_lev5_col44_inst1_port_COUT, FA_lev5_col44_inst2_port_COUT, HA_lev5_col44_inst3_port_COUT, FA_lev4_col45_inst2_port_S, FA_lev4_col45_inst2_port_COUT);
FA_lev4_col46_inst0: FA PORT MAP(FA_lev5_col46_inst0_port_S, FA_lev5_col46_inst1_port_S, HA_lev5_col46_inst2_port_S, FA_lev4_col46_inst0_port_S, FA_lev4_col46_inst0_port_COUT);
FA_lev4_col46_inst1: FA PORT MAP(PP_IN(8)(46), PP_IN(9)(46), PP_IN(10)(46), FA_lev4_col46_inst1_port_S, FA_lev4_col46_inst1_port_COUT);
FA_lev4_col46_inst2: FA PORT MAP(FA_lev5_col45_inst0_port_COUT, FA_lev5_col45_inst1_port_COUT, FA_lev5_col45_inst2_port_COUT, FA_lev4_col46_inst2_port_S, FA_lev4_col46_inst2_port_COUT);
FA_lev4_col47_inst0: FA PORT MAP(FA_lev5_col47_inst0_port_S, FA_lev5_col47_inst1_port_S, PP_IN(6)(47), FA_lev4_col47_inst0_port_S, FA_lev4_col47_inst0_port_COUT);
FA_lev4_col47_inst1: FA PORT MAP(PP_IN(7)(47), PP_IN(8)(47), PP_IN(9)(47), FA_lev4_col47_inst1_port_S, FA_lev4_col47_inst1_port_COUT);
FA_lev4_col47_inst2: FA PORT MAP(FA_lev5_col46_inst0_port_COUT, FA_lev5_col46_inst1_port_COUT, HA_lev5_col46_inst2_port_COUT, FA_lev4_col47_inst2_port_S, FA_lev4_col47_inst2_port_COUT);
FA_lev4_col48_inst0: FA PORT MAP(FA_lev5_col48_inst0_port_S, HA_lev5_col48_inst1_port_S, PP_IN(5)(48), FA_lev4_col48_inst0_port_S, FA_lev4_col48_inst0_port_COUT);
FA_lev4_col48_inst1: FA PORT MAP(PP_IN(6)(48), PP_IN(7)(48), PP_IN(8)(48), FA_lev4_col48_inst1_port_S, FA_lev4_col48_inst1_port_COUT);
FA_lev4_col48_inst2: FA PORT MAP(PP_IN(9)(48), FA_lev5_col47_inst0_port_COUT, FA_lev5_col47_inst1_port_COUT, FA_lev4_col48_inst2_port_S, FA_lev4_col48_inst2_port_COUT);
FA_lev4_col49_inst0: FA PORT MAP(FA_lev5_col49_inst0_port_S, PP_IN(3)(49), PP_IN(4)(49), FA_lev4_col49_inst0_port_S, FA_lev4_col49_inst0_port_COUT);
FA_lev4_col49_inst1: FA PORT MAP(PP_IN(5)(49), PP_IN(6)(49), PP_IN(7)(49), FA_lev4_col49_inst1_port_S, FA_lev4_col49_inst1_port_COUT);
FA_lev4_col49_inst2: FA PORT MAP(PP_IN(8)(49), FA_lev5_col48_inst0_port_COUT, HA_lev5_col48_inst1_port_COUT, FA_lev4_col49_inst2_port_S, FA_lev4_col49_inst2_port_COUT);
FA_lev4_col50_inst0: FA PORT MAP(HA_lev5_col50_inst0_port_S, PP_IN(2)(50), PP_IN(3)(50), FA_lev4_col50_inst0_port_S, FA_lev4_col50_inst0_port_COUT);
FA_lev4_col50_inst1: FA PORT MAP(PP_IN(4)(50), PP_IN(5)(50), PP_IN(6)(50), FA_lev4_col50_inst1_port_S, FA_lev4_col50_inst1_port_COUT);
FA_lev4_col50_inst2: FA PORT MAP(PP_IN(7)(50), PP_IN(8)(50), FA_lev5_col49_inst0_port_COUT, FA_lev4_col50_inst2_port_S, FA_lev4_col50_inst2_port_COUT);
FA_lev4_col51_inst0: FA PORT MAP(PP_IN(0)(51), PP_IN(1)(51), PP_IN(2)(51), FA_lev4_col51_inst0_port_S, FA_lev4_col51_inst0_port_COUT);
FA_lev4_col51_inst1: FA PORT MAP(PP_IN(3)(51), PP_IN(4)(51), PP_IN(5)(51), FA_lev4_col51_inst1_port_S, FA_lev4_col51_inst1_port_COUT);
FA_lev4_col51_inst2: FA PORT MAP(PP_IN(6)(51), PP_IN(7)(51), HA_lev5_col50_inst0_port_COUT, FA_lev4_col51_inst2_port_S, FA_lev4_col51_inst2_port_COUT);
FA_lev4_col52_inst0: FA PORT MAP(PP_IN(0)(52), PP_IN(1)(52), PP_IN(2)(52), FA_lev4_col52_inst0_port_S, FA_lev4_col52_inst0_port_COUT);
FA_lev4_col52_inst1: FA PORT MAP(PP_IN(3)(52), PP_IN(4)(52), PP_IN(5)(52), FA_lev4_col52_inst1_port_S, FA_lev4_col52_inst1_port_COUT);
HA_lev4_col52_inst2: HA PORT MAP(PP_IN(6)(52), PP_IN(7)(52), HA_lev4_col52_inst2_port_S, HA_lev4_col52_inst2_port_COUT);
FA_lev4_col53_inst0: FA PORT MAP(PP_IN(0)(53), PP_IN(1)(53), PP_IN(2)(53), FA_lev4_col53_inst0_port_S, FA_lev4_col53_inst0_port_COUT);
FA_lev4_col53_inst1: FA PORT MAP(PP_IN(3)(53), PP_IN(4)(53), PP_IN(5)(53), FA_lev4_col53_inst1_port_S, FA_lev4_col53_inst1_port_COUT);
FA_lev4_col54_inst0: FA PORT MAP(PP_IN(0)(54), PP_IN(1)(54), PP_IN(2)(54), FA_lev4_col54_inst0_port_S, FA_lev4_col54_inst0_port_COUT);
HA_lev4_col54_inst1: HA PORT MAP(PP_IN(3)(54), PP_IN(4)(54), HA_lev4_col54_inst1_port_S, HA_lev4_col54_inst1_port_COUT);
FA_lev4_col55_inst0: FA PORT MAP(PP_IN(0)(55), PP_IN(1)(55), PP_IN(2)(55), FA_lev4_col55_inst0_port_S, FA_lev4_col55_inst0_port_COUT);
HA_lev4_col56_inst0: HA PORT MAP(PP_IN(0)(56), PP_IN(1)(56), HA_lev4_col56_inst0_port_S, HA_lev4_col56_inst0_port_COUT);

-- Level no 4
HA_lev3_col6_inst0: HA PORT MAP(PP_IN(0)(6), PP_IN(1)(6), HA_lev3_col6_inst0_port_S, HA_lev3_col6_inst0_port_COUT);
HA_lev3_col7_inst0: HA PORT MAP(PP_IN(0)(7), PP_IN(1)(7), HA_lev3_col7_inst0_port_S, HA_lev3_col7_inst0_port_COUT);
FA_lev3_col8_inst0: FA PORT MAP(PP_IN(0)(8), PP_IN(1)(8), PP_IN(2)(8), FA_lev3_col8_inst0_port_S, FA_lev3_col8_inst0_port_COUT);
HA_lev3_col8_inst1: HA PORT MAP(PP_IN(3)(8), PP_IN(4)(8), HA_lev3_col8_inst1_port_S, HA_lev3_col8_inst1_port_COUT);
FA_lev3_col9_inst0: FA PORT MAP(PP_IN(0)(9), PP_IN(1)(9), PP_IN(2)(9), FA_lev3_col9_inst0_port_S, FA_lev3_col9_inst0_port_COUT);
HA_lev3_col9_inst1: HA PORT MAP(PP_IN(3)(9), PP_IN(4)(9), HA_lev3_col9_inst1_port_S, HA_lev3_col9_inst1_port_COUT);
FA_lev3_col10_inst0: FA PORT MAP(HA_lev4_col10_inst0_port_S, PP_IN(2)(10), PP_IN(3)(10), FA_lev3_col10_inst0_port_S, FA_lev3_col10_inst0_port_COUT);
FA_lev3_col10_inst1: FA PORT MAP(PP_IN(4)(10), PP_IN(5)(10), PP_IN(6)(10), FA_lev3_col10_inst1_port_S, FA_lev3_col10_inst1_port_COUT);
FA_lev3_col11_inst0: FA PORT MAP(HA_lev4_col11_inst0_port_S, PP_IN(2)(11), PP_IN(3)(11), FA_lev3_col11_inst0_port_S, FA_lev3_col11_inst0_port_COUT);
FA_lev3_col11_inst1: FA PORT MAP(PP_IN(4)(11), PP_IN(5)(11), HA_lev4_col10_inst0_port_COUT, FA_lev3_col11_inst1_port_S, FA_lev3_col11_inst1_port_COUT);
FA_lev3_col12_inst0: FA PORT MAP(FA_lev4_col12_inst0_port_S, HA_lev4_col12_inst1_port_S, PP_IN(5)(12), FA_lev3_col12_inst0_port_S, FA_lev3_col12_inst0_port_COUT);
FA_lev3_col12_inst1: FA PORT MAP(PP_IN(6)(12), PP_IN(7)(12), HA_lev4_col11_inst0_port_COUT, FA_lev3_col12_inst1_port_S, FA_lev3_col12_inst1_port_COUT);
FA_lev3_col13_inst0: FA PORT MAP(FA_lev4_col13_inst0_port_S, HA_lev4_col13_inst1_port_S, PP_IN(5)(13), FA_lev3_col13_inst0_port_S, FA_lev3_col13_inst0_port_COUT);
FA_lev3_col13_inst1: FA PORT MAP(PP_IN(6)(13), FA_lev4_col12_inst0_port_COUT, HA_lev4_col12_inst1_port_COUT, FA_lev3_col13_inst1_port_S, FA_lev3_col13_inst1_port_COUT);
FA_lev3_col14_inst0: FA PORT MAP(FA_lev4_col14_inst0_port_S, FA_lev4_col14_inst1_port_S, HA_lev4_col14_inst2_port_S, FA_lev3_col14_inst0_port_S, FA_lev3_col14_inst0_port_COUT);
FA_lev3_col14_inst1: FA PORT MAP(PP_IN(8)(14), FA_lev4_col13_inst0_port_COUT, HA_lev4_col13_inst1_port_COUT, FA_lev3_col14_inst1_port_S, FA_lev3_col14_inst1_port_COUT);
FA_lev3_col15_inst0: FA PORT MAP(FA_lev4_col15_inst0_port_S, FA_lev4_col15_inst1_port_S, HA_lev4_col15_inst2_port_S, FA_lev3_col15_inst0_port_S, FA_lev3_col15_inst0_port_COUT);
FA_lev3_col15_inst1: FA PORT MAP(FA_lev4_col14_inst0_port_COUT, FA_lev4_col14_inst1_port_COUT, HA_lev4_col14_inst2_port_COUT, FA_lev3_col15_inst1_port_S, FA_lev3_col15_inst1_port_COUT);
FA_lev3_col16_inst0: FA PORT MAP(FA_lev4_col16_inst0_port_S, FA_lev4_col16_inst1_port_S, FA_lev4_col16_inst2_port_S, FA_lev3_col16_inst0_port_S, FA_lev3_col16_inst0_port_COUT);
FA_lev3_col16_inst1: FA PORT MAP(FA_lev4_col15_inst0_port_COUT, FA_lev4_col15_inst1_port_COUT, HA_lev4_col15_inst2_port_COUT, FA_lev3_col16_inst1_port_S, FA_lev3_col16_inst1_port_COUT);
FA_lev3_col17_inst0: FA PORT MAP(FA_lev4_col17_inst0_port_S, FA_lev4_col17_inst1_port_S, FA_lev4_col17_inst2_port_S, FA_lev3_col17_inst0_port_S, FA_lev3_col17_inst0_port_COUT);
FA_lev3_col17_inst1: FA PORT MAP(FA_lev4_col16_inst0_port_COUT, FA_lev4_col16_inst1_port_COUT, FA_lev4_col16_inst2_port_COUT, FA_lev3_col17_inst1_port_S, FA_lev3_col17_inst1_port_COUT);
FA_lev3_col18_inst0: FA PORT MAP(FA_lev4_col18_inst0_port_S, FA_lev4_col18_inst1_port_S, FA_lev4_col18_inst2_port_S, FA_lev3_col18_inst0_port_S, FA_lev3_col18_inst0_port_COUT);
FA_lev3_col18_inst1: FA PORT MAP(FA_lev4_col17_inst0_port_COUT, FA_lev4_col17_inst1_port_COUT, FA_lev4_col17_inst2_port_COUT, FA_lev3_col18_inst1_port_S, FA_lev3_col18_inst1_port_COUT);
FA_lev3_col19_inst0: FA PORT MAP(FA_lev4_col19_inst0_port_S, FA_lev4_col19_inst1_port_S, FA_lev4_col19_inst2_port_S, FA_lev3_col19_inst0_port_S, FA_lev3_col19_inst0_port_COUT);
FA_lev3_col19_inst1: FA PORT MAP(FA_lev4_col18_inst0_port_COUT, FA_lev4_col18_inst1_port_COUT, FA_lev4_col18_inst2_port_COUT, FA_lev3_col19_inst1_port_S, FA_lev3_col19_inst1_port_COUT);
FA_lev3_col20_inst0: FA PORT MAP(FA_lev4_col20_inst0_port_S, FA_lev4_col20_inst1_port_S, FA_lev4_col20_inst2_port_S, FA_lev3_col20_inst0_port_S, FA_lev3_col20_inst0_port_COUT);
FA_lev3_col20_inst1: FA PORT MAP(FA_lev4_col19_inst0_port_COUT, FA_lev4_col19_inst1_port_COUT, FA_lev4_col19_inst2_port_COUT, FA_lev3_col20_inst1_port_S, FA_lev3_col20_inst1_port_COUT);
FA_lev3_col21_inst0: FA PORT MAP(FA_lev4_col21_inst0_port_S, FA_lev4_col21_inst1_port_S, FA_lev4_col21_inst2_port_S, FA_lev3_col21_inst0_port_S, FA_lev3_col21_inst0_port_COUT);
FA_lev3_col21_inst1: FA PORT MAP(FA_lev4_col20_inst0_port_COUT, FA_lev4_col20_inst1_port_COUT, FA_lev4_col20_inst2_port_COUT, FA_lev3_col21_inst1_port_S, FA_lev3_col21_inst1_port_COUT);
FA_lev3_col22_inst0: FA PORT MAP(FA_lev4_col22_inst0_port_S, FA_lev4_col22_inst1_port_S, FA_lev4_col22_inst2_port_S, FA_lev3_col22_inst0_port_S, FA_lev3_col22_inst0_port_COUT);
FA_lev3_col22_inst1: FA PORT MAP(FA_lev4_col21_inst0_port_COUT, FA_lev4_col21_inst1_port_COUT, FA_lev4_col21_inst2_port_COUT, FA_lev3_col22_inst1_port_S, FA_lev3_col22_inst1_port_COUT);
FA_lev3_col23_inst0: FA PORT MAP(FA_lev4_col23_inst0_port_S, FA_lev4_col23_inst1_port_S, FA_lev4_col23_inst2_port_S, FA_lev3_col23_inst0_port_S, FA_lev3_col23_inst0_port_COUT);
FA_lev3_col23_inst1: FA PORT MAP(FA_lev4_col22_inst0_port_COUT, FA_lev4_col22_inst1_port_COUT, FA_lev4_col22_inst2_port_COUT, FA_lev3_col23_inst1_port_S, FA_lev3_col23_inst1_port_COUT);
FA_lev3_col24_inst0: FA PORT MAP(FA_lev4_col24_inst0_port_S, FA_lev4_col24_inst1_port_S, FA_lev4_col24_inst2_port_S, FA_lev3_col24_inst0_port_S, FA_lev3_col24_inst0_port_COUT);
FA_lev3_col24_inst1: FA PORT MAP(FA_lev4_col23_inst0_port_COUT, FA_lev4_col23_inst1_port_COUT, FA_lev4_col23_inst2_port_COUT, FA_lev3_col24_inst1_port_S, FA_lev3_col24_inst1_port_COUT);
FA_lev3_col25_inst0: FA PORT MAP(FA_lev4_col25_inst0_port_S, FA_lev4_col25_inst1_port_S, FA_lev4_col25_inst2_port_S, FA_lev3_col25_inst0_port_S, FA_lev3_col25_inst0_port_COUT);
FA_lev3_col25_inst1: FA PORT MAP(FA_lev4_col24_inst0_port_COUT, FA_lev4_col24_inst1_port_COUT, FA_lev4_col24_inst2_port_COUT, FA_lev3_col25_inst1_port_S, FA_lev3_col25_inst1_port_COUT);
FA_lev3_col26_inst0: FA PORT MAP(FA_lev4_col26_inst0_port_S, FA_lev4_col26_inst1_port_S, FA_lev4_col26_inst2_port_S, FA_lev3_col26_inst0_port_S, FA_lev3_col26_inst0_port_COUT);
FA_lev3_col26_inst1: FA PORT MAP(FA_lev4_col25_inst0_port_COUT, FA_lev4_col25_inst1_port_COUT, FA_lev4_col25_inst2_port_COUT, FA_lev3_col26_inst1_port_S, FA_lev3_col26_inst1_port_COUT);
FA_lev3_col27_inst0: FA PORT MAP(FA_lev4_col27_inst0_port_S, FA_lev4_col27_inst1_port_S, FA_lev4_col27_inst2_port_S, FA_lev3_col27_inst0_port_S, FA_lev3_col27_inst0_port_COUT);
FA_lev3_col27_inst1: FA PORT MAP(FA_lev4_col26_inst0_port_COUT, FA_lev4_col26_inst1_port_COUT, FA_lev4_col26_inst2_port_COUT, FA_lev3_col27_inst1_port_S, FA_lev3_col27_inst1_port_COUT);
FA_lev3_col28_inst0: FA PORT MAP(FA_lev4_col28_inst0_port_S, FA_lev4_col28_inst1_port_S, FA_lev4_col28_inst2_port_S, FA_lev3_col28_inst0_port_S, FA_lev3_col28_inst0_port_COUT);
FA_lev3_col28_inst1: FA PORT MAP(FA_lev4_col27_inst0_port_COUT, FA_lev4_col27_inst1_port_COUT, FA_lev4_col27_inst2_port_COUT, FA_lev3_col28_inst1_port_S, FA_lev3_col28_inst1_port_COUT);
FA_lev3_col29_inst0: FA PORT MAP(FA_lev4_col29_inst0_port_S, FA_lev4_col29_inst1_port_S, FA_lev4_col29_inst2_port_S, FA_lev3_col29_inst0_port_S, FA_lev3_col29_inst0_port_COUT);
FA_lev3_col29_inst1: FA PORT MAP(FA_lev4_col28_inst0_port_COUT, FA_lev4_col28_inst1_port_COUT, FA_lev4_col28_inst2_port_COUT, FA_lev3_col29_inst1_port_S, FA_lev3_col29_inst1_port_COUT);
FA_lev3_col30_inst0: FA PORT MAP(FA_lev4_col30_inst0_port_S, FA_lev4_col30_inst1_port_S, FA_lev4_col30_inst2_port_S, FA_lev3_col30_inst0_port_S, FA_lev3_col30_inst0_port_COUT);
FA_lev3_col30_inst1: FA PORT MAP(FA_lev4_col29_inst0_port_COUT, FA_lev4_col29_inst1_port_COUT, FA_lev4_col29_inst2_port_COUT, FA_lev3_col30_inst1_port_S, FA_lev3_col30_inst1_port_COUT);
FA_lev3_col31_inst0: FA PORT MAP(FA_lev4_col31_inst0_port_S, FA_lev4_col31_inst1_port_S, FA_lev4_col31_inst2_port_S, FA_lev3_col31_inst0_port_S, FA_lev3_col31_inst0_port_COUT);
FA_lev3_col31_inst1: FA PORT MAP(FA_lev4_col30_inst0_port_COUT, FA_lev4_col30_inst1_port_COUT, FA_lev4_col30_inst2_port_COUT, FA_lev3_col31_inst1_port_S, FA_lev3_col31_inst1_port_COUT);
FA_lev3_col32_inst0: FA PORT MAP(FA_lev4_col32_inst0_port_S, FA_lev4_col32_inst1_port_S, FA_lev4_col32_inst2_port_S, FA_lev3_col32_inst0_port_S, FA_lev3_col32_inst0_port_COUT);
FA_lev3_col32_inst1: FA PORT MAP(FA_lev4_col31_inst0_port_COUT, FA_lev4_col31_inst1_port_COUT, FA_lev4_col31_inst2_port_COUT, FA_lev3_col32_inst1_port_S, FA_lev3_col32_inst1_port_COUT);
FA_lev3_col33_inst0: FA PORT MAP(FA_lev4_col33_inst0_port_S, FA_lev4_col33_inst1_port_S, FA_lev4_col33_inst2_port_S, FA_lev3_col33_inst0_port_S, FA_lev3_col33_inst0_port_COUT);
FA_lev3_col33_inst1: FA PORT MAP(FA_lev4_col32_inst0_port_COUT, FA_lev4_col32_inst1_port_COUT, FA_lev4_col32_inst2_port_COUT, FA_lev3_col33_inst1_port_S, FA_lev3_col33_inst1_port_COUT);
FA_lev3_col34_inst0: FA PORT MAP(FA_lev4_col34_inst0_port_S, FA_lev4_col34_inst1_port_S, FA_lev4_col34_inst2_port_S, FA_lev3_col34_inst0_port_S, FA_lev3_col34_inst0_port_COUT);
FA_lev3_col34_inst1: FA PORT MAP(FA_lev4_col33_inst0_port_COUT, FA_lev4_col33_inst1_port_COUT, FA_lev4_col33_inst2_port_COUT, FA_lev3_col34_inst1_port_S, FA_lev3_col34_inst1_port_COUT);
FA_lev3_col35_inst0: FA PORT MAP(FA_lev4_col35_inst0_port_S, FA_lev4_col35_inst1_port_S, FA_lev4_col35_inst2_port_S, FA_lev3_col35_inst0_port_S, FA_lev3_col35_inst0_port_COUT);
FA_lev3_col35_inst1: FA PORT MAP(FA_lev4_col34_inst0_port_COUT, FA_lev4_col34_inst1_port_COUT, FA_lev4_col34_inst2_port_COUT, FA_lev3_col35_inst1_port_S, FA_lev3_col35_inst1_port_COUT);
FA_lev3_col36_inst0: FA PORT MAP(FA_lev4_col36_inst0_port_S, FA_lev4_col36_inst1_port_S, FA_lev4_col36_inst2_port_S, FA_lev3_col36_inst0_port_S, FA_lev3_col36_inst0_port_COUT);
FA_lev3_col36_inst1: FA PORT MAP(FA_lev4_col35_inst0_port_COUT, FA_lev4_col35_inst1_port_COUT, FA_lev4_col35_inst2_port_COUT, FA_lev3_col36_inst1_port_S, FA_lev3_col36_inst1_port_COUT);
FA_lev3_col37_inst0: FA PORT MAP(FA_lev4_col37_inst0_port_S, FA_lev4_col37_inst1_port_S, FA_lev4_col37_inst2_port_S, FA_lev3_col37_inst0_port_S, FA_lev3_col37_inst0_port_COUT);
FA_lev3_col37_inst1: FA PORT MAP(FA_lev4_col36_inst0_port_COUT, FA_lev4_col36_inst1_port_COUT, FA_lev4_col36_inst2_port_COUT, FA_lev3_col37_inst1_port_S, FA_lev3_col37_inst1_port_COUT);
FA_lev3_col38_inst0: FA PORT MAP(FA_lev4_col38_inst0_port_S, FA_lev4_col38_inst1_port_S, FA_lev4_col38_inst2_port_S, FA_lev3_col38_inst0_port_S, FA_lev3_col38_inst0_port_COUT);
FA_lev3_col38_inst1: FA PORT MAP(FA_lev4_col37_inst0_port_COUT, FA_lev4_col37_inst1_port_COUT, FA_lev4_col37_inst2_port_COUT, FA_lev3_col38_inst1_port_S, FA_lev3_col38_inst1_port_COUT);
FA_lev3_col39_inst0: FA PORT MAP(FA_lev4_col39_inst0_port_S, FA_lev4_col39_inst1_port_S, FA_lev4_col39_inst2_port_S, FA_lev3_col39_inst0_port_S, FA_lev3_col39_inst0_port_COUT);
FA_lev3_col39_inst1: FA PORT MAP(FA_lev4_col38_inst0_port_COUT, FA_lev4_col38_inst1_port_COUT, FA_lev4_col38_inst2_port_COUT, FA_lev3_col39_inst1_port_S, FA_lev3_col39_inst1_port_COUT);
FA_lev3_col40_inst0: FA PORT MAP(FA_lev4_col40_inst0_port_S, FA_lev4_col40_inst1_port_S, FA_lev4_col40_inst2_port_S, FA_lev3_col40_inst0_port_S, FA_lev3_col40_inst0_port_COUT);
FA_lev3_col40_inst1: FA PORT MAP(FA_lev4_col39_inst0_port_COUT, FA_lev4_col39_inst1_port_COUT, FA_lev4_col39_inst2_port_COUT, FA_lev3_col40_inst1_port_S, FA_lev3_col40_inst1_port_COUT);
FA_lev3_col41_inst0: FA PORT MAP(FA_lev4_col41_inst0_port_S, FA_lev4_col41_inst1_port_S, FA_lev4_col41_inst2_port_S, FA_lev3_col41_inst0_port_S, FA_lev3_col41_inst0_port_COUT);
FA_lev3_col41_inst1: FA PORT MAP(FA_lev4_col40_inst0_port_COUT, FA_lev4_col40_inst1_port_COUT, FA_lev4_col40_inst2_port_COUT, FA_lev3_col41_inst1_port_S, FA_lev3_col41_inst1_port_COUT);
FA_lev3_col42_inst0: FA PORT MAP(FA_lev4_col42_inst0_port_S, FA_lev4_col42_inst1_port_S, FA_lev4_col42_inst2_port_S, FA_lev3_col42_inst0_port_S, FA_lev3_col42_inst0_port_COUT);
FA_lev3_col42_inst1: FA PORT MAP(FA_lev4_col41_inst0_port_COUT, FA_lev4_col41_inst1_port_COUT, FA_lev4_col41_inst2_port_COUT, FA_lev3_col42_inst1_port_S, FA_lev3_col42_inst1_port_COUT);
FA_lev3_col43_inst0: FA PORT MAP(FA_lev4_col43_inst0_port_S, FA_lev4_col43_inst1_port_S, FA_lev4_col43_inst2_port_S, FA_lev3_col43_inst0_port_S, FA_lev3_col43_inst0_port_COUT);
FA_lev3_col43_inst1: FA PORT MAP(FA_lev4_col42_inst0_port_COUT, FA_lev4_col42_inst1_port_COUT, FA_lev4_col42_inst2_port_COUT, FA_lev3_col43_inst1_port_S, FA_lev3_col43_inst1_port_COUT);
FA_lev3_col44_inst0: FA PORT MAP(FA_lev4_col44_inst0_port_S, FA_lev4_col44_inst1_port_S, FA_lev4_col44_inst2_port_S, FA_lev3_col44_inst0_port_S, FA_lev3_col44_inst0_port_COUT);
FA_lev3_col44_inst1: FA PORT MAP(FA_lev4_col43_inst0_port_COUT, FA_lev4_col43_inst1_port_COUT, FA_lev4_col43_inst2_port_COUT, FA_lev3_col44_inst1_port_S, FA_lev3_col44_inst1_port_COUT);
FA_lev3_col45_inst0: FA PORT MAP(FA_lev4_col45_inst0_port_S, FA_lev4_col45_inst1_port_S, FA_lev4_col45_inst2_port_S, FA_lev3_col45_inst0_port_S, FA_lev3_col45_inst0_port_COUT);
FA_lev3_col45_inst1: FA PORT MAP(FA_lev4_col44_inst0_port_COUT, FA_lev4_col44_inst1_port_COUT, FA_lev4_col44_inst2_port_COUT, FA_lev3_col45_inst1_port_S, FA_lev3_col45_inst1_port_COUT);
FA_lev3_col46_inst0: FA PORT MAP(FA_lev4_col46_inst0_port_S, FA_lev4_col46_inst1_port_S, FA_lev4_col46_inst2_port_S, FA_lev3_col46_inst0_port_S, FA_lev3_col46_inst0_port_COUT);
FA_lev3_col46_inst1: FA PORT MAP(FA_lev4_col45_inst0_port_COUT, FA_lev4_col45_inst1_port_COUT, FA_lev4_col45_inst2_port_COUT, FA_lev3_col46_inst1_port_S, FA_lev3_col46_inst1_port_COUT);
FA_lev3_col47_inst0: FA PORT MAP(FA_lev4_col47_inst0_port_S, FA_lev4_col47_inst1_port_S, FA_lev4_col47_inst2_port_S, FA_lev3_col47_inst0_port_S, FA_lev3_col47_inst0_port_COUT);
FA_lev3_col47_inst1: FA PORT MAP(FA_lev4_col46_inst0_port_COUT, FA_lev4_col46_inst1_port_COUT, FA_lev4_col46_inst2_port_COUT, FA_lev3_col47_inst1_port_S, FA_lev3_col47_inst1_port_COUT);
FA_lev3_col48_inst0: FA PORT MAP(FA_lev4_col48_inst0_port_S, FA_lev4_col48_inst1_port_S, FA_lev4_col48_inst2_port_S, FA_lev3_col48_inst0_port_S, FA_lev3_col48_inst0_port_COUT);
FA_lev3_col48_inst1: FA PORT MAP(FA_lev4_col47_inst0_port_COUT, FA_lev4_col47_inst1_port_COUT, FA_lev4_col47_inst2_port_COUT, FA_lev3_col48_inst1_port_S, FA_lev3_col48_inst1_port_COUT);
FA_lev3_col49_inst0: FA PORT MAP(FA_lev4_col49_inst0_port_S, FA_lev4_col49_inst1_port_S, FA_lev4_col49_inst2_port_S, FA_lev3_col49_inst0_port_S, FA_lev3_col49_inst0_port_COUT);
FA_lev3_col49_inst1: FA PORT MAP(FA_lev4_col48_inst0_port_COUT, FA_lev4_col48_inst1_port_COUT, FA_lev4_col48_inst2_port_COUT, FA_lev3_col49_inst1_port_S, FA_lev3_col49_inst1_port_COUT);
FA_lev3_col50_inst0: FA PORT MAP(FA_lev4_col50_inst0_port_S, FA_lev4_col50_inst1_port_S, FA_lev4_col50_inst2_port_S, FA_lev3_col50_inst0_port_S, FA_lev3_col50_inst0_port_COUT);
FA_lev3_col50_inst1: FA PORT MAP(FA_lev4_col49_inst0_port_COUT, FA_lev4_col49_inst1_port_COUT, FA_lev4_col49_inst2_port_COUT, FA_lev3_col50_inst1_port_S, FA_lev3_col50_inst1_port_COUT);
FA_lev3_col51_inst0: FA PORT MAP(FA_lev4_col51_inst0_port_S, FA_lev4_col51_inst1_port_S, FA_lev4_col51_inst2_port_S, FA_lev3_col51_inst0_port_S, FA_lev3_col51_inst0_port_COUT);
FA_lev3_col51_inst1: FA PORT MAP(FA_lev4_col50_inst0_port_COUT, FA_lev4_col50_inst1_port_COUT, FA_lev4_col50_inst2_port_COUT, FA_lev3_col51_inst1_port_S, FA_lev3_col51_inst1_port_COUT);
FA_lev3_col52_inst0: FA PORT MAP(FA_lev4_col52_inst0_port_S, FA_lev4_col52_inst1_port_S, HA_lev4_col52_inst2_port_S, FA_lev3_col52_inst0_port_S, FA_lev3_col52_inst0_port_COUT);
FA_lev3_col52_inst1: FA PORT MAP(FA_lev4_col51_inst0_port_COUT, FA_lev4_col51_inst1_port_COUT, FA_lev4_col51_inst2_port_COUT, FA_lev3_col52_inst1_port_S, FA_lev3_col52_inst1_port_COUT);
FA_lev3_col53_inst0: FA PORT MAP(FA_lev4_col53_inst0_port_S, FA_lev4_col53_inst1_port_S, PP_IN(6)(53), FA_lev3_col53_inst0_port_S, FA_lev3_col53_inst0_port_COUT);
FA_lev3_col53_inst1: FA PORT MAP(FA_lev4_col52_inst0_port_COUT, FA_lev4_col52_inst1_port_COUT, HA_lev4_col52_inst2_port_COUT, FA_lev3_col53_inst1_port_S, FA_lev3_col53_inst1_port_COUT);
FA_lev3_col54_inst0: FA PORT MAP(FA_lev4_col54_inst0_port_S, HA_lev4_col54_inst1_port_S, PP_IN(5)(54), FA_lev3_col54_inst0_port_S, FA_lev3_col54_inst0_port_COUT);
FA_lev3_col54_inst1: FA PORT MAP(PP_IN(6)(54), FA_lev4_col53_inst0_port_COUT, FA_lev4_col53_inst1_port_COUT, FA_lev3_col54_inst1_port_S, FA_lev3_col54_inst1_port_COUT);
FA_lev3_col55_inst0: FA PORT MAP(FA_lev4_col55_inst0_port_S, PP_IN(3)(55), PP_IN(4)(55), FA_lev3_col55_inst0_port_S, FA_lev3_col55_inst0_port_COUT);
FA_lev3_col55_inst1: FA PORT MAP(PP_IN(5)(55), FA_lev4_col54_inst0_port_COUT, HA_lev4_col54_inst1_port_COUT, FA_lev3_col55_inst1_port_S, FA_lev3_col55_inst1_port_COUT);
FA_lev3_col56_inst0: FA PORT MAP(HA_lev4_col56_inst0_port_S, PP_IN(2)(56), PP_IN(3)(56), FA_lev3_col56_inst0_port_S, FA_lev3_col56_inst0_port_COUT);
FA_lev3_col56_inst1: FA PORT MAP(PP_IN(4)(56), PP_IN(5)(56), FA_lev4_col55_inst0_port_COUT, FA_lev3_col56_inst1_port_S, FA_lev3_col56_inst1_port_COUT);
FA_lev3_col57_inst0: FA PORT MAP(PP_IN(0)(57), PP_IN(1)(57), PP_IN(2)(57), FA_lev3_col57_inst0_port_S, FA_lev3_col57_inst0_port_COUT);
FA_lev3_col57_inst1: FA PORT MAP(PP_IN(3)(57), PP_IN(4)(57), HA_lev4_col56_inst0_port_COUT, FA_lev3_col57_inst1_port_S, FA_lev3_col57_inst1_port_COUT);
FA_lev3_col58_inst0: FA PORT MAP(PP_IN(0)(58), PP_IN(1)(58), PP_IN(2)(58), FA_lev3_col58_inst0_port_S, FA_lev3_col58_inst0_port_COUT);
HA_lev3_col58_inst1: HA PORT MAP(PP_IN(3)(58), PP_IN(4)(58), HA_lev3_col58_inst1_port_S, HA_lev3_col58_inst1_port_COUT);
FA_lev3_col59_inst0: FA PORT MAP(PP_IN(0)(59), PP_IN(1)(59), PP_IN(2)(59), FA_lev3_col59_inst0_port_S, FA_lev3_col59_inst0_port_COUT);
HA_lev3_col60_inst0: HA PORT MAP(PP_IN(0)(60), PP_IN(1)(60), HA_lev3_col60_inst0_port_S, HA_lev3_col60_inst0_port_COUT);

-- Level no 3
HA_lev2_col4_inst0: HA PORT MAP(PP_IN(0)(4), PP_IN(1)(4), HA_lev2_col4_inst0_port_S, HA_lev2_col4_inst0_port_COUT);
HA_lev2_col5_inst0: HA PORT MAP(PP_IN(0)(5), PP_IN(1)(5), HA_lev2_col5_inst0_port_S, HA_lev2_col5_inst0_port_COUT);
FA_lev2_col6_inst0: FA PORT MAP(HA_lev3_col6_inst0_port_S, PP_IN(2)(6), PP_IN(3)(6), FA_lev2_col6_inst0_port_S, FA_lev2_col6_inst0_port_COUT);
FA_lev2_col7_inst0: FA PORT MAP(HA_lev3_col7_inst0_port_S, PP_IN(2)(7), PP_IN(3)(7), FA_lev2_col7_inst0_port_S, FA_lev2_col7_inst0_port_COUT);
FA_lev2_col8_inst0: FA PORT MAP(FA_lev3_col8_inst0_port_S, HA_lev3_col8_inst1_port_S, PP_IN(5)(8), FA_lev2_col8_inst0_port_S, FA_lev2_col8_inst0_port_COUT);
FA_lev2_col9_inst0: FA PORT MAP(FA_lev3_col9_inst0_port_S, HA_lev3_col9_inst1_port_S, FA_lev3_col8_inst0_port_COUT, FA_lev2_col9_inst0_port_S, FA_lev2_col9_inst0_port_COUT);
FA_lev2_col10_inst0: FA PORT MAP(FA_lev3_col10_inst0_port_S, FA_lev3_col10_inst1_port_S, FA_lev3_col9_inst0_port_COUT, FA_lev2_col10_inst0_port_S, FA_lev2_col10_inst0_port_COUT);
FA_lev2_col11_inst0: FA PORT MAP(FA_lev3_col11_inst0_port_S, FA_lev3_col11_inst1_port_S, FA_lev3_col10_inst0_port_COUT, FA_lev2_col11_inst0_port_S, FA_lev2_col11_inst0_port_COUT);
FA_lev2_col12_inst0: FA PORT MAP(FA_lev3_col12_inst0_port_S, FA_lev3_col12_inst1_port_S, FA_lev3_col11_inst0_port_COUT, FA_lev2_col12_inst0_port_S, FA_lev2_col12_inst0_port_COUT);
FA_lev2_col13_inst0: FA PORT MAP(FA_lev3_col13_inst0_port_S, FA_lev3_col13_inst1_port_S, FA_lev3_col12_inst0_port_COUT, FA_lev2_col13_inst0_port_S, FA_lev2_col13_inst0_port_COUT);
FA_lev2_col14_inst0: FA PORT MAP(FA_lev3_col14_inst0_port_S, FA_lev3_col14_inst1_port_S, FA_lev3_col13_inst0_port_COUT, FA_lev2_col14_inst0_port_S, FA_lev2_col14_inst0_port_COUT);
FA_lev2_col15_inst0: FA PORT MAP(FA_lev3_col15_inst0_port_S, FA_lev3_col15_inst1_port_S, FA_lev3_col14_inst0_port_COUT, FA_lev2_col15_inst0_port_S, FA_lev2_col15_inst0_port_COUT);
FA_lev2_col16_inst0: FA PORT MAP(FA_lev3_col16_inst0_port_S, FA_lev3_col16_inst1_port_S, FA_lev3_col15_inst0_port_COUT, FA_lev2_col16_inst0_port_S, FA_lev2_col16_inst0_port_COUT);
FA_lev2_col17_inst0: FA PORT MAP(FA_lev3_col17_inst0_port_S, FA_lev3_col17_inst1_port_S, FA_lev3_col16_inst0_port_COUT, FA_lev2_col17_inst0_port_S, FA_lev2_col17_inst0_port_COUT);
FA_lev2_col18_inst0: FA PORT MAP(FA_lev3_col18_inst0_port_S, FA_lev3_col18_inst1_port_S, FA_lev3_col17_inst0_port_COUT, FA_lev2_col18_inst0_port_S, FA_lev2_col18_inst0_port_COUT);
FA_lev2_col19_inst0: FA PORT MAP(FA_lev3_col19_inst0_port_S, FA_lev3_col19_inst1_port_S, FA_lev3_col18_inst0_port_COUT, FA_lev2_col19_inst0_port_S, FA_lev2_col19_inst0_port_COUT);
FA_lev2_col20_inst0: FA PORT MAP(FA_lev3_col20_inst0_port_S, FA_lev3_col20_inst1_port_S, FA_lev3_col19_inst0_port_COUT, FA_lev2_col20_inst0_port_S, FA_lev2_col20_inst0_port_COUT);
FA_lev2_col21_inst0: FA PORT MAP(FA_lev3_col21_inst0_port_S, FA_lev3_col21_inst1_port_S, FA_lev3_col20_inst0_port_COUT, FA_lev2_col21_inst0_port_S, FA_lev2_col21_inst0_port_COUT);
FA_lev2_col22_inst0: FA PORT MAP(FA_lev3_col22_inst0_port_S, FA_lev3_col22_inst1_port_S, FA_lev3_col21_inst0_port_COUT, FA_lev2_col22_inst0_port_S, FA_lev2_col22_inst0_port_COUT);
FA_lev2_col23_inst0: FA PORT MAP(FA_lev3_col23_inst0_port_S, FA_lev3_col23_inst1_port_S, FA_lev3_col22_inst0_port_COUT, FA_lev2_col23_inst0_port_S, FA_lev2_col23_inst0_port_COUT);
FA_lev2_col24_inst0: FA PORT MAP(FA_lev3_col24_inst0_port_S, FA_lev3_col24_inst1_port_S, FA_lev3_col23_inst0_port_COUT, FA_lev2_col24_inst0_port_S, FA_lev2_col24_inst0_port_COUT);
FA_lev2_col25_inst0: FA PORT MAP(FA_lev3_col25_inst0_port_S, FA_lev3_col25_inst1_port_S, FA_lev3_col24_inst0_port_COUT, FA_lev2_col25_inst0_port_S, FA_lev2_col25_inst0_port_COUT);
FA_lev2_col26_inst0: FA PORT MAP(FA_lev3_col26_inst0_port_S, FA_lev3_col26_inst1_port_S, FA_lev3_col25_inst0_port_COUT, FA_lev2_col26_inst0_port_S, FA_lev2_col26_inst0_port_COUT);
FA_lev2_col27_inst0: FA PORT MAP(FA_lev3_col27_inst0_port_S, FA_lev3_col27_inst1_port_S, FA_lev3_col26_inst0_port_COUT, FA_lev2_col27_inst0_port_S, FA_lev2_col27_inst0_port_COUT);
FA_lev2_col28_inst0: FA PORT MAP(FA_lev3_col28_inst0_port_S, FA_lev3_col28_inst1_port_S, FA_lev3_col27_inst0_port_COUT, FA_lev2_col28_inst0_port_S, FA_lev2_col28_inst0_port_COUT);
FA_lev2_col29_inst0: FA PORT MAP(FA_lev3_col29_inst0_port_S, FA_lev3_col29_inst1_port_S, FA_lev3_col28_inst0_port_COUT, FA_lev2_col29_inst0_port_S, FA_lev2_col29_inst0_port_COUT);
FA_lev2_col30_inst0: FA PORT MAP(FA_lev3_col30_inst0_port_S, FA_lev3_col30_inst1_port_S, FA_lev3_col29_inst0_port_COUT, FA_lev2_col30_inst0_port_S, FA_lev2_col30_inst0_port_COUT);
FA_lev2_col31_inst0: FA PORT MAP(FA_lev3_col31_inst0_port_S, FA_lev3_col31_inst1_port_S, FA_lev3_col30_inst0_port_COUT, FA_lev2_col31_inst0_port_S, FA_lev2_col31_inst0_port_COUT);
FA_lev2_col32_inst0: FA PORT MAP(FA_lev3_col32_inst0_port_S, FA_lev3_col32_inst1_port_S, FA_lev3_col31_inst0_port_COUT, FA_lev2_col32_inst0_port_S, FA_lev2_col32_inst0_port_COUT);
FA_lev2_col33_inst0: FA PORT MAP(FA_lev3_col33_inst0_port_S, FA_lev3_col33_inst1_port_S, FA_lev3_col32_inst0_port_COUT, FA_lev2_col33_inst0_port_S, FA_lev2_col33_inst0_port_COUT);
FA_lev2_col34_inst0: FA PORT MAP(FA_lev3_col34_inst0_port_S, FA_lev3_col34_inst1_port_S, FA_lev3_col33_inst0_port_COUT, FA_lev2_col34_inst0_port_S, FA_lev2_col34_inst0_port_COUT);
FA_lev2_col35_inst0: FA PORT MAP(FA_lev3_col35_inst0_port_S, FA_lev3_col35_inst1_port_S, FA_lev3_col34_inst0_port_COUT, FA_lev2_col35_inst0_port_S, FA_lev2_col35_inst0_port_COUT);
FA_lev2_col36_inst0: FA PORT MAP(FA_lev3_col36_inst0_port_S, FA_lev3_col36_inst1_port_S, FA_lev3_col35_inst0_port_COUT, FA_lev2_col36_inst0_port_S, FA_lev2_col36_inst0_port_COUT);
FA_lev2_col37_inst0: FA PORT MAP(FA_lev3_col37_inst0_port_S, FA_lev3_col37_inst1_port_S, FA_lev3_col36_inst0_port_COUT, FA_lev2_col37_inst0_port_S, FA_lev2_col37_inst0_port_COUT);
FA_lev2_col38_inst0: FA PORT MAP(FA_lev3_col38_inst0_port_S, FA_lev3_col38_inst1_port_S, FA_lev3_col37_inst0_port_COUT, FA_lev2_col38_inst0_port_S, FA_lev2_col38_inst0_port_COUT);
FA_lev2_col39_inst0: FA PORT MAP(FA_lev3_col39_inst0_port_S, FA_lev3_col39_inst1_port_S, FA_lev3_col38_inst0_port_COUT, FA_lev2_col39_inst0_port_S, FA_lev2_col39_inst0_port_COUT);
FA_lev2_col40_inst0: FA PORT MAP(FA_lev3_col40_inst0_port_S, FA_lev3_col40_inst1_port_S, FA_lev3_col39_inst0_port_COUT, FA_lev2_col40_inst0_port_S, FA_lev2_col40_inst0_port_COUT);
FA_lev2_col41_inst0: FA PORT MAP(FA_lev3_col41_inst0_port_S, FA_lev3_col41_inst1_port_S, FA_lev3_col40_inst0_port_COUT, FA_lev2_col41_inst0_port_S, FA_lev2_col41_inst0_port_COUT);
FA_lev2_col42_inst0: FA PORT MAP(FA_lev3_col42_inst0_port_S, FA_lev3_col42_inst1_port_S, FA_lev3_col41_inst0_port_COUT, FA_lev2_col42_inst0_port_S, FA_lev2_col42_inst0_port_COUT);
FA_lev2_col43_inst0: FA PORT MAP(FA_lev3_col43_inst0_port_S, FA_lev3_col43_inst1_port_S, FA_lev3_col42_inst0_port_COUT, FA_lev2_col43_inst0_port_S, FA_lev2_col43_inst0_port_COUT);
FA_lev2_col44_inst0: FA PORT MAP(FA_lev3_col44_inst0_port_S, FA_lev3_col44_inst1_port_S, FA_lev3_col43_inst0_port_COUT, FA_lev2_col44_inst0_port_S, FA_lev2_col44_inst0_port_COUT);
FA_lev2_col45_inst0: FA PORT MAP(FA_lev3_col45_inst0_port_S, FA_lev3_col45_inst1_port_S, FA_lev3_col44_inst0_port_COUT, FA_lev2_col45_inst0_port_S, FA_lev2_col45_inst0_port_COUT);
FA_lev2_col46_inst0: FA PORT MAP(FA_lev3_col46_inst0_port_S, FA_lev3_col46_inst1_port_S, FA_lev3_col45_inst0_port_COUT, FA_lev2_col46_inst0_port_S, FA_lev2_col46_inst0_port_COUT);
FA_lev2_col47_inst0: FA PORT MAP(FA_lev3_col47_inst0_port_S, FA_lev3_col47_inst1_port_S, FA_lev3_col46_inst0_port_COUT, FA_lev2_col47_inst0_port_S, FA_lev2_col47_inst0_port_COUT);
FA_lev2_col48_inst0: FA PORT MAP(FA_lev3_col48_inst0_port_S, FA_lev3_col48_inst1_port_S, FA_lev3_col47_inst0_port_COUT, FA_lev2_col48_inst0_port_S, FA_lev2_col48_inst0_port_COUT);
FA_lev2_col49_inst0: FA PORT MAP(FA_lev3_col49_inst0_port_S, FA_lev3_col49_inst1_port_S, FA_lev3_col48_inst0_port_COUT, FA_lev2_col49_inst0_port_S, FA_lev2_col49_inst0_port_COUT);
FA_lev2_col50_inst0: FA PORT MAP(FA_lev3_col50_inst0_port_S, FA_lev3_col50_inst1_port_S, FA_lev3_col49_inst0_port_COUT, FA_lev2_col50_inst0_port_S, FA_lev2_col50_inst0_port_COUT);
FA_lev2_col51_inst0: FA PORT MAP(FA_lev3_col51_inst0_port_S, FA_lev3_col51_inst1_port_S, FA_lev3_col50_inst0_port_COUT, FA_lev2_col51_inst0_port_S, FA_lev2_col51_inst0_port_COUT);
FA_lev2_col52_inst0: FA PORT MAP(FA_lev3_col52_inst0_port_S, FA_lev3_col52_inst1_port_S, FA_lev3_col51_inst0_port_COUT, FA_lev2_col52_inst0_port_S, FA_lev2_col52_inst0_port_COUT);
FA_lev2_col53_inst0: FA PORT MAP(FA_lev3_col53_inst0_port_S, FA_lev3_col53_inst1_port_S, FA_lev3_col52_inst0_port_COUT, FA_lev2_col53_inst0_port_S, FA_lev2_col53_inst0_port_COUT);
FA_lev2_col54_inst0: FA PORT MAP(FA_lev3_col54_inst0_port_S, FA_lev3_col54_inst1_port_S, FA_lev3_col53_inst0_port_COUT, FA_lev2_col54_inst0_port_S, FA_lev2_col54_inst0_port_COUT);
FA_lev2_col55_inst0: FA PORT MAP(FA_lev3_col55_inst0_port_S, FA_lev3_col55_inst1_port_S, FA_lev3_col54_inst0_port_COUT, FA_lev2_col55_inst0_port_S, FA_lev2_col55_inst0_port_COUT);
FA_lev2_col56_inst0: FA PORT MAP(FA_lev3_col56_inst0_port_S, FA_lev3_col56_inst1_port_S, FA_lev3_col55_inst0_port_COUT, FA_lev2_col56_inst0_port_S, FA_lev2_col56_inst0_port_COUT);
FA_lev2_col57_inst0: FA PORT MAP(FA_lev3_col57_inst0_port_S, FA_lev3_col57_inst1_port_S, FA_lev3_col56_inst0_port_COUT, FA_lev2_col57_inst0_port_S, FA_lev2_col57_inst0_port_COUT);
FA_lev2_col58_inst0: FA PORT MAP(FA_lev3_col58_inst0_port_S, HA_lev3_col58_inst1_port_S, FA_lev3_col57_inst0_port_COUT, FA_lev2_col58_inst0_port_S, FA_lev2_col58_inst0_port_COUT);
FA_lev2_col59_inst0: FA PORT MAP(FA_lev3_col59_inst0_port_S, PP_IN(3)(59), FA_lev3_col58_inst0_port_COUT, FA_lev2_col59_inst0_port_S, FA_lev2_col59_inst0_port_COUT);
FA_lev2_col60_inst0: FA PORT MAP(HA_lev3_col60_inst0_port_S, PP_IN(2)(60), PP_IN(3)(60), FA_lev2_col60_inst0_port_S, FA_lev2_col60_inst0_port_COUT);
FA_lev2_col61_inst0: FA PORT MAP(PP_IN(0)(61), PP_IN(1)(61), PP_IN(2)(61), FA_lev2_col61_inst0_port_S, FA_lev2_col61_inst0_port_COUT);
HA_lev2_col62_inst0: HA PORT MAP(PP_IN(0)(62), PP_IN(1)(62), HA_lev2_col62_inst0_port_S, HA_lev2_col62_inst0_port_COUT);

-- Level no 2
HA_lev1_col2_inst0: HA PORT MAP(PP_IN(0)(2), PP_IN(1)(2), HA_lev1_col2_inst0_port_S, HA_lev1_col2_inst0_port_COUT);
HA_lev1_col3_inst0: HA PORT MAP(PP_IN(0)(3), PP_IN(1)(3), HA_lev1_col3_inst0_port_S, HA_lev1_col3_inst0_port_COUT);
FA_lev1_col4_inst0: FA PORT MAP(HA_lev2_col4_inst0_port_S, PP_IN(2)(4), PP_IN(3)(4), FA_lev1_col4_inst0_port_S, FA_lev1_col4_inst0_port_COUT);
FA_lev1_col5_inst0: FA PORT MAP(HA_lev2_col5_inst0_port_S, PP_IN(2)(5), HA_lev2_col4_inst0_port_COUT, FA_lev1_col5_inst0_port_S, FA_lev1_col5_inst0_port_COUT);
FA_lev1_col6_inst0: FA PORT MAP(FA_lev2_col6_inst0_port_S, PP_IN(4)(6), HA_lev2_col5_inst0_port_COUT, FA_lev1_col6_inst0_port_S, FA_lev1_col6_inst0_port_COUT);
FA_lev1_col7_inst0: FA PORT MAP(FA_lev2_col7_inst0_port_S, HA_lev3_col6_inst0_port_COUT, FA_lev2_col6_inst0_port_COUT, FA_lev1_col7_inst0_port_S, FA_lev1_col7_inst0_port_COUT);
FA_lev1_col8_inst0: FA PORT MAP(FA_lev2_col8_inst0_port_S, HA_lev3_col7_inst0_port_COUT, FA_lev2_col7_inst0_port_COUT, FA_lev1_col8_inst0_port_S, FA_lev1_col8_inst0_port_COUT);
FA_lev1_col9_inst0: FA PORT MAP(FA_lev2_col9_inst0_port_S, HA_lev3_col8_inst1_port_COUT, FA_lev2_col8_inst0_port_COUT, FA_lev1_col9_inst0_port_S, FA_lev1_col9_inst0_port_COUT);
FA_lev1_col10_inst0: FA PORT MAP(FA_lev2_col10_inst0_port_S, HA_lev3_col9_inst1_port_COUT, FA_lev2_col9_inst0_port_COUT, FA_lev1_col10_inst0_port_S, FA_lev1_col10_inst0_port_COUT);
FA_lev1_col11_inst0: FA PORT MAP(FA_lev2_col11_inst0_port_S, FA_lev3_col10_inst1_port_COUT, FA_lev2_col10_inst0_port_COUT, FA_lev1_col11_inst0_port_S, FA_lev1_col11_inst0_port_COUT);
FA_lev1_col12_inst0: FA PORT MAP(FA_lev2_col12_inst0_port_S, FA_lev3_col11_inst1_port_COUT, FA_lev2_col11_inst0_port_COUT, FA_lev1_col12_inst0_port_S, FA_lev1_col12_inst0_port_COUT);
FA_lev1_col13_inst0: FA PORT MAP(FA_lev2_col13_inst0_port_S, FA_lev3_col12_inst1_port_COUT, FA_lev2_col12_inst0_port_COUT, FA_lev1_col13_inst0_port_S, FA_lev1_col13_inst0_port_COUT);
FA_lev1_col14_inst0: FA PORT MAP(FA_lev2_col14_inst0_port_S, FA_lev3_col13_inst1_port_COUT, FA_lev2_col13_inst0_port_COUT, FA_lev1_col14_inst0_port_S, FA_lev1_col14_inst0_port_COUT);
FA_lev1_col15_inst0: FA PORT MAP(FA_lev2_col15_inst0_port_S, FA_lev3_col14_inst1_port_COUT, FA_lev2_col14_inst0_port_COUT, FA_lev1_col15_inst0_port_S, FA_lev1_col15_inst0_port_COUT);
FA_lev1_col16_inst0: FA PORT MAP(FA_lev2_col16_inst0_port_S, FA_lev3_col15_inst1_port_COUT, FA_lev2_col15_inst0_port_COUT, FA_lev1_col16_inst0_port_S, FA_lev1_col16_inst0_port_COUT);
FA_lev1_col17_inst0: FA PORT MAP(FA_lev2_col17_inst0_port_S, FA_lev3_col16_inst1_port_COUT, FA_lev2_col16_inst0_port_COUT, FA_lev1_col17_inst0_port_S, FA_lev1_col17_inst0_port_COUT);
FA_lev1_col18_inst0: FA PORT MAP(FA_lev2_col18_inst0_port_S, FA_lev3_col17_inst1_port_COUT, FA_lev2_col17_inst0_port_COUT, FA_lev1_col18_inst0_port_S, FA_lev1_col18_inst0_port_COUT);
FA_lev1_col19_inst0: FA PORT MAP(FA_lev2_col19_inst0_port_S, FA_lev3_col18_inst1_port_COUT, FA_lev2_col18_inst0_port_COUT, FA_lev1_col19_inst0_port_S, FA_lev1_col19_inst0_port_COUT);
FA_lev1_col20_inst0: FA PORT MAP(FA_lev2_col20_inst0_port_S, FA_lev3_col19_inst1_port_COUT, FA_lev2_col19_inst0_port_COUT, FA_lev1_col20_inst0_port_S, FA_lev1_col20_inst0_port_COUT);
FA_lev1_col21_inst0: FA PORT MAP(FA_lev2_col21_inst0_port_S, FA_lev3_col20_inst1_port_COUT, FA_lev2_col20_inst0_port_COUT, FA_lev1_col21_inst0_port_S, FA_lev1_col21_inst0_port_COUT);
FA_lev1_col22_inst0: FA PORT MAP(FA_lev2_col22_inst0_port_S, FA_lev3_col21_inst1_port_COUT, FA_lev2_col21_inst0_port_COUT, FA_lev1_col22_inst0_port_S, FA_lev1_col22_inst0_port_COUT);
FA_lev1_col23_inst0: FA PORT MAP(FA_lev2_col23_inst0_port_S, FA_lev3_col22_inst1_port_COUT, FA_lev2_col22_inst0_port_COUT, FA_lev1_col23_inst0_port_S, FA_lev1_col23_inst0_port_COUT);
FA_lev1_col24_inst0: FA PORT MAP(FA_lev2_col24_inst0_port_S, FA_lev3_col23_inst1_port_COUT, FA_lev2_col23_inst0_port_COUT, FA_lev1_col24_inst0_port_S, FA_lev1_col24_inst0_port_COUT);
FA_lev1_col25_inst0: FA PORT MAP(FA_lev2_col25_inst0_port_S, FA_lev3_col24_inst1_port_COUT, FA_lev2_col24_inst0_port_COUT, FA_lev1_col25_inst0_port_S, FA_lev1_col25_inst0_port_COUT);
FA_lev1_col26_inst0: FA PORT MAP(FA_lev2_col26_inst0_port_S, FA_lev3_col25_inst1_port_COUT, FA_lev2_col25_inst0_port_COUT, FA_lev1_col26_inst0_port_S, FA_lev1_col26_inst0_port_COUT);
FA_lev1_col27_inst0: FA PORT MAP(FA_lev2_col27_inst0_port_S, FA_lev3_col26_inst1_port_COUT, FA_lev2_col26_inst0_port_COUT, FA_lev1_col27_inst0_port_S, FA_lev1_col27_inst0_port_COUT);
FA_lev1_col28_inst0: FA PORT MAP(FA_lev2_col28_inst0_port_S, FA_lev3_col27_inst1_port_COUT, FA_lev2_col27_inst0_port_COUT, FA_lev1_col28_inst0_port_S, FA_lev1_col28_inst0_port_COUT);
FA_lev1_col29_inst0: FA PORT MAP(FA_lev2_col29_inst0_port_S, FA_lev3_col28_inst1_port_COUT, FA_lev2_col28_inst0_port_COUT, FA_lev1_col29_inst0_port_S, FA_lev1_col29_inst0_port_COUT);
FA_lev1_col30_inst0: FA PORT MAP(FA_lev2_col30_inst0_port_S, FA_lev3_col29_inst1_port_COUT, FA_lev2_col29_inst0_port_COUT, FA_lev1_col30_inst0_port_S, FA_lev1_col30_inst0_port_COUT);
FA_lev1_col31_inst0: FA PORT MAP(FA_lev2_col31_inst0_port_S, FA_lev3_col30_inst1_port_COUT, FA_lev2_col30_inst0_port_COUT, FA_lev1_col31_inst0_port_S, FA_lev1_col31_inst0_port_COUT);
FA_lev1_col32_inst0: FA PORT MAP(FA_lev2_col32_inst0_port_S, FA_lev3_col31_inst1_port_COUT, FA_lev2_col31_inst0_port_COUT, FA_lev1_col32_inst0_port_S, FA_lev1_col32_inst0_port_COUT);
FA_lev1_col33_inst0: FA PORT MAP(FA_lev2_col33_inst0_port_S, FA_lev3_col32_inst1_port_COUT, FA_lev2_col32_inst0_port_COUT, FA_lev1_col33_inst0_port_S, FA_lev1_col33_inst0_port_COUT);
FA_lev1_col34_inst0: FA PORT MAP(FA_lev2_col34_inst0_port_S, FA_lev3_col33_inst1_port_COUT, FA_lev2_col33_inst0_port_COUT, FA_lev1_col34_inst0_port_S, FA_lev1_col34_inst0_port_COUT);
FA_lev1_col35_inst0: FA PORT MAP(FA_lev2_col35_inst0_port_S, FA_lev3_col34_inst1_port_COUT, FA_lev2_col34_inst0_port_COUT, FA_lev1_col35_inst0_port_S, FA_lev1_col35_inst0_port_COUT);
FA_lev1_col36_inst0: FA PORT MAP(FA_lev2_col36_inst0_port_S, FA_lev3_col35_inst1_port_COUT, FA_lev2_col35_inst0_port_COUT, FA_lev1_col36_inst0_port_S, FA_lev1_col36_inst0_port_COUT);
FA_lev1_col37_inst0: FA PORT MAP(FA_lev2_col37_inst0_port_S, FA_lev3_col36_inst1_port_COUT, FA_lev2_col36_inst0_port_COUT, FA_lev1_col37_inst0_port_S, FA_lev1_col37_inst0_port_COUT);
FA_lev1_col38_inst0: FA PORT MAP(FA_lev2_col38_inst0_port_S, FA_lev3_col37_inst1_port_COUT, FA_lev2_col37_inst0_port_COUT, FA_lev1_col38_inst0_port_S, FA_lev1_col38_inst0_port_COUT);
FA_lev1_col39_inst0: FA PORT MAP(FA_lev2_col39_inst0_port_S, FA_lev3_col38_inst1_port_COUT, FA_lev2_col38_inst0_port_COUT, FA_lev1_col39_inst0_port_S, FA_lev1_col39_inst0_port_COUT);
FA_lev1_col40_inst0: FA PORT MAP(FA_lev2_col40_inst0_port_S, FA_lev3_col39_inst1_port_COUT, FA_lev2_col39_inst0_port_COUT, FA_lev1_col40_inst0_port_S, FA_lev1_col40_inst0_port_COUT);
FA_lev1_col41_inst0: FA PORT MAP(FA_lev2_col41_inst0_port_S, FA_lev3_col40_inst1_port_COUT, FA_lev2_col40_inst0_port_COUT, FA_lev1_col41_inst0_port_S, FA_lev1_col41_inst0_port_COUT);
FA_lev1_col42_inst0: FA PORT MAP(FA_lev2_col42_inst0_port_S, FA_lev3_col41_inst1_port_COUT, FA_lev2_col41_inst0_port_COUT, FA_lev1_col42_inst0_port_S, FA_lev1_col42_inst0_port_COUT);
FA_lev1_col43_inst0: FA PORT MAP(FA_lev2_col43_inst0_port_S, FA_lev3_col42_inst1_port_COUT, FA_lev2_col42_inst0_port_COUT, FA_lev1_col43_inst0_port_S, FA_lev1_col43_inst0_port_COUT);
FA_lev1_col44_inst0: FA PORT MAP(FA_lev2_col44_inst0_port_S, FA_lev3_col43_inst1_port_COUT, FA_lev2_col43_inst0_port_COUT, FA_lev1_col44_inst0_port_S, FA_lev1_col44_inst0_port_COUT);
FA_lev1_col45_inst0: FA PORT MAP(FA_lev2_col45_inst0_port_S, FA_lev3_col44_inst1_port_COUT, FA_lev2_col44_inst0_port_COUT, FA_lev1_col45_inst0_port_S, FA_lev1_col45_inst0_port_COUT);
FA_lev1_col46_inst0: FA PORT MAP(FA_lev2_col46_inst0_port_S, FA_lev3_col45_inst1_port_COUT, FA_lev2_col45_inst0_port_COUT, FA_lev1_col46_inst0_port_S, FA_lev1_col46_inst0_port_COUT);
FA_lev1_col47_inst0: FA PORT MAP(FA_lev2_col47_inst0_port_S, FA_lev3_col46_inst1_port_COUT, FA_lev2_col46_inst0_port_COUT, FA_lev1_col47_inst0_port_S, FA_lev1_col47_inst0_port_COUT);
FA_lev1_col48_inst0: FA PORT MAP(FA_lev2_col48_inst0_port_S, FA_lev3_col47_inst1_port_COUT, FA_lev2_col47_inst0_port_COUT, FA_lev1_col48_inst0_port_S, FA_lev1_col48_inst0_port_COUT);
FA_lev1_col49_inst0: FA PORT MAP(FA_lev2_col49_inst0_port_S, FA_lev3_col48_inst1_port_COUT, FA_lev2_col48_inst0_port_COUT, FA_lev1_col49_inst0_port_S, FA_lev1_col49_inst0_port_COUT);
FA_lev1_col50_inst0: FA PORT MAP(FA_lev2_col50_inst0_port_S, FA_lev3_col49_inst1_port_COUT, FA_lev2_col49_inst0_port_COUT, FA_lev1_col50_inst0_port_S, FA_lev1_col50_inst0_port_COUT);
FA_lev1_col51_inst0: FA PORT MAP(FA_lev2_col51_inst0_port_S, FA_lev3_col50_inst1_port_COUT, FA_lev2_col50_inst0_port_COUT, FA_lev1_col51_inst0_port_S, FA_lev1_col51_inst0_port_COUT);
FA_lev1_col52_inst0: FA PORT MAP(FA_lev2_col52_inst0_port_S, FA_lev3_col51_inst1_port_COUT, FA_lev2_col51_inst0_port_COUT, FA_lev1_col52_inst0_port_S, FA_lev1_col52_inst0_port_COUT);
FA_lev1_col53_inst0: FA PORT MAP(FA_lev2_col53_inst0_port_S, FA_lev3_col52_inst1_port_COUT, FA_lev2_col52_inst0_port_COUT, FA_lev1_col53_inst0_port_S, FA_lev1_col53_inst0_port_COUT);
FA_lev1_col54_inst0: FA PORT MAP(FA_lev2_col54_inst0_port_S, FA_lev3_col53_inst1_port_COUT, FA_lev2_col53_inst0_port_COUT, FA_lev1_col54_inst0_port_S, FA_lev1_col54_inst0_port_COUT);
FA_lev1_col55_inst0: FA PORT MAP(FA_lev2_col55_inst0_port_S, FA_lev3_col54_inst1_port_COUT, FA_lev2_col54_inst0_port_COUT, FA_lev1_col55_inst0_port_S, FA_lev1_col55_inst0_port_COUT);
FA_lev1_col56_inst0: FA PORT MAP(FA_lev2_col56_inst0_port_S, FA_lev3_col55_inst1_port_COUT, FA_lev2_col55_inst0_port_COUT, FA_lev1_col56_inst0_port_S, FA_lev1_col56_inst0_port_COUT);
FA_lev1_col57_inst0: FA PORT MAP(FA_lev2_col57_inst0_port_S, FA_lev3_col56_inst1_port_COUT, FA_lev2_col56_inst0_port_COUT, FA_lev1_col57_inst0_port_S, FA_lev1_col57_inst0_port_COUT);
FA_lev1_col58_inst0: FA PORT MAP(FA_lev2_col58_inst0_port_S, FA_lev3_col57_inst1_port_COUT, FA_lev2_col57_inst0_port_COUT, FA_lev1_col58_inst0_port_S, FA_lev1_col58_inst0_port_COUT);
FA_lev1_col59_inst0: FA PORT MAP(FA_lev2_col59_inst0_port_S, HA_lev3_col58_inst1_port_COUT, FA_lev2_col58_inst0_port_COUT, FA_lev1_col59_inst0_port_S, FA_lev1_col59_inst0_port_COUT);
FA_lev1_col60_inst0: FA PORT MAP(FA_lev2_col60_inst0_port_S, FA_lev3_col59_inst0_port_COUT, FA_lev2_col59_inst0_port_COUT, FA_lev1_col60_inst0_port_S, FA_lev1_col60_inst0_port_COUT);
FA_lev1_col61_inst0: FA PORT MAP(FA_lev2_col61_inst0_port_S, HA_lev3_col60_inst0_port_COUT, FA_lev2_col60_inst0_port_COUT, FA_lev1_col61_inst0_port_S, FA_lev1_col61_inst0_port_COUT);
FA_lev1_col62_inst0: FA PORT MAP(HA_lev2_col62_inst0_port_S, PP_IN(2)(62), FA_lev2_col61_inst0_port_COUT, FA_lev1_col62_inst0_port_S, FA_lev1_col62_inst0_port_COUT);
FA_lev1_col63_inst0: FA PORT MAP(PP_IN(0)(63), PP_IN(1)(63), HA_lev2_col62_inst0_port_COUT, FA_lev1_col63_inst0_port_S, FA_lev1_col63_inst0_port_COUT);


PP_OUT1 <=  FA_lev1_col63_inst0_port_S & FA_lev1_col62_inst0_port_S & FA_lev1_col61_inst0_port_S & FA_lev1_col60_inst0_port_S & FA_lev1_col59_inst0_port_S & FA_lev1_col58_inst0_port_S & FA_lev1_col57_inst0_port_S & FA_lev1_col56_inst0_port_S & FA_lev1_col55_inst0_port_S & FA_lev1_col54_inst0_port_S & FA_lev1_col53_inst0_port_S & FA_lev1_col52_inst0_port_S & FA_lev1_col51_inst0_port_S & FA_lev1_col50_inst0_port_S & FA_lev1_col49_inst0_port_S & FA_lev1_col48_inst0_port_S & FA_lev1_col47_inst0_port_S & FA_lev1_col46_inst0_port_S & FA_lev1_col45_inst0_port_S & FA_lev1_col44_inst0_port_S & FA_lev1_col43_inst0_port_S & FA_lev1_col42_inst0_port_S & FA_lev1_col41_inst0_port_S & FA_lev1_col40_inst0_port_S & FA_lev1_col39_inst0_port_S & FA_lev1_col38_inst0_port_S & FA_lev1_col37_inst0_port_S & FA_lev1_col36_inst0_port_S & FA_lev1_col35_inst0_port_S & FA_lev1_col34_inst0_port_S & FA_lev1_col33_inst0_port_S & FA_lev1_col32_inst0_port_S & FA_lev1_col31_inst0_port_S & FA_lev1_col30_inst0_port_S & FA_lev1_col29_inst0_port_S & FA_lev1_col28_inst0_port_S & FA_lev1_col27_inst0_port_S & FA_lev1_col26_inst0_port_S & FA_lev1_col25_inst0_port_S & FA_lev1_col24_inst0_port_S & FA_lev1_col23_inst0_port_S & FA_lev1_col22_inst0_port_S & FA_lev1_col21_inst0_port_S & FA_lev1_col20_inst0_port_S & FA_lev1_col19_inst0_port_S & FA_lev1_col18_inst0_port_S & FA_lev1_col17_inst0_port_S & FA_lev1_col16_inst0_port_S & FA_lev1_col15_inst0_port_S & FA_lev1_col14_inst0_port_S & FA_lev1_col13_inst0_port_S & FA_lev1_col12_inst0_port_S & FA_lev1_col11_inst0_port_S & FA_lev1_col10_inst0_port_S & FA_lev1_col9_inst0_port_S & FA_lev1_col8_inst0_port_S & FA_lev1_col7_inst0_port_S & FA_lev1_col6_inst0_port_S & FA_lev1_col5_inst0_port_S & FA_lev1_col4_inst0_port_S & HA_lev1_col3_inst0_port_S & HA_lev1_col2_inst0_port_S & PP_IN(0)(1) & PP_IN(0)(0);

PP_OUT2 <=  FA_lev1_col62_inst0_port_COUT & FA_lev1_col61_inst0_port_COUT & FA_lev1_col60_inst0_port_COUT & FA_lev1_col59_inst0_port_COUT & FA_lev1_col58_inst0_port_COUT & FA_lev1_col57_inst0_port_COUT & FA_lev1_col56_inst0_port_COUT & FA_lev1_col55_inst0_port_COUT & FA_lev1_col54_inst0_port_COUT & FA_lev1_col53_inst0_port_COUT & FA_lev1_col52_inst0_port_COUT & FA_lev1_col51_inst0_port_COUT & FA_lev1_col50_inst0_port_COUT & FA_lev1_col49_inst0_port_COUT & FA_lev1_col48_inst0_port_COUT & FA_lev1_col47_inst0_port_COUT & FA_lev1_col46_inst0_port_COUT & FA_lev1_col45_inst0_port_COUT & FA_lev1_col44_inst0_port_COUT & FA_lev1_col43_inst0_port_COUT & FA_lev1_col42_inst0_port_COUT & FA_lev1_col41_inst0_port_COUT & FA_lev1_col40_inst0_port_COUT & FA_lev1_col39_inst0_port_COUT & FA_lev1_col38_inst0_port_COUT & FA_lev1_col37_inst0_port_COUT & FA_lev1_col36_inst0_port_COUT & FA_lev1_col35_inst0_port_COUT & FA_lev1_col34_inst0_port_COUT & FA_lev1_col33_inst0_port_COUT & FA_lev1_col32_inst0_port_COUT & FA_lev1_col31_inst0_port_COUT & FA_lev1_col30_inst0_port_COUT & FA_lev1_col29_inst0_port_COUT & FA_lev1_col28_inst0_port_COUT & FA_lev1_col27_inst0_port_COUT & FA_lev1_col26_inst0_port_COUT & FA_lev1_col25_inst0_port_COUT & FA_lev1_col24_inst0_port_COUT & FA_lev1_col23_inst0_port_COUT & FA_lev1_col22_inst0_port_COUT & FA_lev1_col21_inst0_port_COUT & FA_lev1_col20_inst0_port_COUT & FA_lev1_col19_inst0_port_COUT & FA_lev1_col18_inst0_port_COUT & FA_lev1_col17_inst0_port_COUT & FA_lev1_col16_inst0_port_COUT & FA_lev1_col15_inst0_port_COUT & FA_lev1_col14_inst0_port_COUT & FA_lev1_col13_inst0_port_COUT & FA_lev1_col12_inst0_port_COUT & FA_lev1_col11_inst0_port_COUT & FA_lev1_col10_inst0_port_COUT & FA_lev1_col9_inst0_port_COUT & FA_lev1_col8_inst0_port_COUT & FA_lev1_col7_inst0_port_COUT & FA_lev1_col6_inst0_port_COUT & FA_lev1_col5_inst0_port_COUT & FA_lev1_col4_inst0_port_COUT & HA_lev1_col3_inst0_port_COUT & HA_lev1_col2_inst0_port_COUT & PP_IN(2)(2) & '0' & PP_IN(1)(0);

END ARCHITECTURE;