`ifndef MY_DEFINES
	`define MY_DEFINES
		parameter nb=10;
`endif
